
module cache ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N30, N31, N32, n4179, \CACHE[7][153] , \CACHE[7][149] ,
         \CACHE[7][148] , \CACHE[7][143] , \CACHE[7][142] , \CACHE[7][141] ,
         \CACHE[7][139] , \CACHE[7][138] , \CACHE[7][137] , \CACHE[7][136] ,
         \CACHE[7][132] , \CACHE[7][131] , \CACHE[7][129] , \CACHE[7][128] ,
         \CACHE[7][127] , \CACHE[7][126] , \CACHE[7][125] , \CACHE[7][124] ,
         \CACHE[7][123] , \CACHE[7][122] , \CACHE[7][121] , \CACHE[7][120] ,
         \CACHE[7][119] , \CACHE[7][118] , \CACHE[7][117] , \CACHE[7][116] ,
         \CACHE[7][115] , \CACHE[7][114] , \CACHE[7][113] , \CACHE[7][112] ,
         \CACHE[7][111] , \CACHE[7][110] , \CACHE[7][109] , \CACHE[7][108] ,
         \CACHE[7][107] , \CACHE[7][106] , \CACHE[7][105] , \CACHE[7][104] ,
         \CACHE[7][103] , \CACHE[7][102] , \CACHE[7][101] , \CACHE[7][100] ,
         \CACHE[7][99] , \CACHE[7][98] , \CACHE[7][97] , \CACHE[7][96] ,
         \CACHE[7][95] , \CACHE[7][94] , \CACHE[7][93] , \CACHE[7][92] ,
         \CACHE[7][91] , \CACHE[7][90] , \CACHE[7][89] , \CACHE[7][88] ,
         \CACHE[7][87] , \CACHE[7][86] , \CACHE[7][85] , \CACHE[7][84] ,
         \CACHE[7][83] , \CACHE[7][82] , \CACHE[7][81] , \CACHE[7][80] ,
         \CACHE[7][79] , \CACHE[7][78] , \CACHE[7][77] , \CACHE[7][76] ,
         \CACHE[7][75] , \CACHE[7][74] , \CACHE[7][73] , \CACHE[7][72] ,
         \CACHE[7][71] , \CACHE[7][70] , \CACHE[7][69] , \CACHE[7][68] ,
         \CACHE[7][67] , \CACHE[7][66] , \CACHE[7][65] , \CACHE[7][64] ,
         \CACHE[7][63] , \CACHE[7][62] , \CACHE[7][61] , \CACHE[7][60] ,
         \CACHE[7][59] , \CACHE[7][58] , \CACHE[7][57] , \CACHE[7][56] ,
         \CACHE[7][55] , \CACHE[7][54] , \CACHE[7][53] , \CACHE[7][52] ,
         \CACHE[7][51] , \CACHE[7][50] , \CACHE[7][49] , \CACHE[7][48] ,
         \CACHE[7][47] , \CACHE[7][46] , \CACHE[7][45] , \CACHE[7][44] ,
         \CACHE[7][43] , \CACHE[7][42] , \CACHE[7][41] , \CACHE[7][40] ,
         \CACHE[7][39] , \CACHE[7][38] , \CACHE[7][37] , \CACHE[7][36] ,
         \CACHE[7][35] , \CACHE[7][34] , \CACHE[7][33] , \CACHE[7][32] ,
         \CACHE[7][31] , \CACHE[7][30] , \CACHE[7][29] , \CACHE[7][28] ,
         \CACHE[7][27] , \CACHE[7][26] , \CACHE[7][25] , \CACHE[7][24] ,
         \CACHE[7][23] , \CACHE[7][22] , \CACHE[7][21] , \CACHE[7][20] ,
         \CACHE[7][19] , \CACHE[7][18] , \CACHE[7][17] , \CACHE[7][16] ,
         \CACHE[7][15] , \CACHE[7][14] , \CACHE[7][13] , \CACHE[7][12] ,
         \CACHE[7][11] , \CACHE[7][10] , \CACHE[7][9] , \CACHE[7][8] ,
         \CACHE[7][7] , \CACHE[7][6] , \CACHE[7][5] , \CACHE[7][4] ,
         \CACHE[7][3] , \CACHE[7][2] , \CACHE[7][1] , \CACHE[7][0] ,
         \CACHE[6][153] , \CACHE[6][149] , \CACHE[6][148] , \CACHE[6][143] ,
         \CACHE[6][142] , \CACHE[6][141] , \CACHE[6][139] , \CACHE[6][138] ,
         \CACHE[6][137] , \CACHE[6][136] , \CACHE[6][132] , \CACHE[6][131] ,
         \CACHE[6][129] , \CACHE[6][128] , \CACHE[6][127] , \CACHE[6][126] ,
         \CACHE[6][125] , \CACHE[6][124] , \CACHE[6][123] , \CACHE[6][122] ,
         \CACHE[6][121] , \CACHE[6][120] , \CACHE[6][119] , \CACHE[6][118] ,
         \CACHE[6][117] , \CACHE[6][116] , \CACHE[6][115] , \CACHE[6][114] ,
         \CACHE[6][113] , \CACHE[6][112] , \CACHE[6][111] , \CACHE[6][110] ,
         \CACHE[6][109] , \CACHE[6][108] , \CACHE[6][107] , \CACHE[6][106] ,
         \CACHE[6][105] , \CACHE[6][104] , \CACHE[6][103] , \CACHE[6][102] ,
         \CACHE[6][101] , \CACHE[6][100] , \CACHE[6][99] , \CACHE[6][98] ,
         \CACHE[6][97] , \CACHE[6][96] , \CACHE[6][95] , \CACHE[6][94] ,
         \CACHE[6][93] , \CACHE[6][92] , \CACHE[6][91] , \CACHE[6][90] ,
         \CACHE[6][89] , \CACHE[6][88] , \CACHE[6][87] , \CACHE[6][86] ,
         \CACHE[6][85] , \CACHE[6][84] , \CACHE[6][83] , \CACHE[6][82] ,
         \CACHE[6][81] , \CACHE[6][80] , \CACHE[6][79] , \CACHE[6][78] ,
         \CACHE[6][77] , \CACHE[6][76] , \CACHE[6][75] , \CACHE[6][74] ,
         \CACHE[6][73] , \CACHE[6][72] , \CACHE[6][71] , \CACHE[6][70] ,
         \CACHE[6][69] , \CACHE[6][68] , \CACHE[6][67] , \CACHE[6][66] ,
         \CACHE[6][65] , \CACHE[6][64] , \CACHE[6][63] , \CACHE[6][62] ,
         \CACHE[6][61] , \CACHE[6][60] , \CACHE[6][59] , \CACHE[6][58] ,
         \CACHE[6][57] , \CACHE[6][56] , \CACHE[6][55] , \CACHE[6][54] ,
         \CACHE[6][53] , \CACHE[6][52] , \CACHE[6][51] , \CACHE[6][50] ,
         \CACHE[6][49] , \CACHE[6][48] , \CACHE[6][47] , \CACHE[6][46] ,
         \CACHE[6][45] , \CACHE[6][44] , \CACHE[6][43] , \CACHE[6][42] ,
         \CACHE[6][41] , \CACHE[6][40] , \CACHE[6][39] , \CACHE[6][38] ,
         \CACHE[6][37] , \CACHE[6][36] , \CACHE[6][35] , \CACHE[6][34] ,
         \CACHE[6][33] , \CACHE[6][32] , \CACHE[6][31] , \CACHE[6][30] ,
         \CACHE[6][29] , \CACHE[6][28] , \CACHE[6][27] , \CACHE[6][26] ,
         \CACHE[6][25] , \CACHE[6][24] , \CACHE[6][23] , \CACHE[6][22] ,
         \CACHE[6][21] , \CACHE[6][20] , \CACHE[6][19] , \CACHE[6][18] ,
         \CACHE[6][17] , \CACHE[6][16] , \CACHE[6][15] , \CACHE[6][14] ,
         \CACHE[6][13] , \CACHE[6][12] , \CACHE[6][11] , \CACHE[6][10] ,
         \CACHE[6][9] , \CACHE[6][8] , \CACHE[6][7] , \CACHE[6][6] ,
         \CACHE[6][5] , \CACHE[6][4] , \CACHE[6][3] , \CACHE[6][2] ,
         \CACHE[6][1] , \CACHE[6][0] , \CACHE[5][153] , \CACHE[5][149] ,
         \CACHE[5][148] , \CACHE[5][143] , \CACHE[5][142] , \CACHE[5][141] ,
         \CACHE[5][139] , \CACHE[5][138] , \CACHE[5][137] , \CACHE[5][136] ,
         \CACHE[5][132] , \CACHE[5][131] , \CACHE[5][129] , \CACHE[5][128] ,
         \CACHE[5][127] , \CACHE[5][126] , \CACHE[5][125] , \CACHE[5][124] ,
         \CACHE[5][123] , \CACHE[5][122] , \CACHE[5][121] , \CACHE[5][120] ,
         \CACHE[5][119] , \CACHE[5][118] , \CACHE[5][117] , \CACHE[5][116] ,
         \CACHE[5][115] , \CACHE[5][114] , \CACHE[5][113] , \CACHE[5][112] ,
         \CACHE[5][111] , \CACHE[5][110] , \CACHE[5][109] , \CACHE[5][108] ,
         \CACHE[5][107] , \CACHE[5][106] , \CACHE[5][105] , \CACHE[5][104] ,
         \CACHE[5][103] , \CACHE[5][102] , \CACHE[5][101] , \CACHE[5][100] ,
         \CACHE[5][99] , \CACHE[5][98] , \CACHE[5][97] , \CACHE[5][96] ,
         \CACHE[5][95] , \CACHE[5][94] , \CACHE[5][93] , \CACHE[5][92] ,
         \CACHE[5][91] , \CACHE[5][90] , \CACHE[5][89] , \CACHE[5][88] ,
         \CACHE[5][87] , \CACHE[5][86] , \CACHE[5][85] , \CACHE[5][84] ,
         \CACHE[5][83] , \CACHE[5][82] , \CACHE[5][81] , \CACHE[5][80] ,
         \CACHE[5][79] , \CACHE[5][78] , \CACHE[5][77] , \CACHE[5][76] ,
         \CACHE[5][75] , \CACHE[5][74] , \CACHE[5][73] , \CACHE[5][72] ,
         \CACHE[5][71] , \CACHE[5][70] , \CACHE[5][69] , \CACHE[5][68] ,
         \CACHE[5][67] , \CACHE[5][66] , \CACHE[5][65] , \CACHE[5][64] ,
         \CACHE[5][63] , \CACHE[5][62] , \CACHE[5][61] , \CACHE[5][60] ,
         \CACHE[5][59] , \CACHE[5][58] , \CACHE[5][57] , \CACHE[5][56] ,
         \CACHE[5][55] , \CACHE[5][54] , \CACHE[5][53] , \CACHE[5][52] ,
         \CACHE[5][51] , \CACHE[5][50] , \CACHE[5][49] , \CACHE[5][48] ,
         \CACHE[5][47] , \CACHE[5][46] , \CACHE[5][45] , \CACHE[5][44] ,
         \CACHE[5][43] , \CACHE[5][42] , \CACHE[5][41] , \CACHE[5][40] ,
         \CACHE[5][39] , \CACHE[5][38] , \CACHE[5][37] , \CACHE[5][36] ,
         \CACHE[5][35] , \CACHE[5][34] , \CACHE[5][33] , \CACHE[5][32] ,
         \CACHE[5][31] , \CACHE[5][30] , \CACHE[5][29] , \CACHE[5][28] ,
         \CACHE[5][27] , \CACHE[5][26] , \CACHE[5][25] , \CACHE[5][24] ,
         \CACHE[5][23] , \CACHE[5][22] , \CACHE[5][21] , \CACHE[5][20] ,
         \CACHE[5][19] , \CACHE[5][18] , \CACHE[5][17] , \CACHE[5][16] ,
         \CACHE[5][15] , \CACHE[5][14] , \CACHE[5][13] , \CACHE[5][12] ,
         \CACHE[5][11] , \CACHE[5][10] , \CACHE[5][9] , \CACHE[5][8] ,
         \CACHE[5][7] , \CACHE[5][6] , \CACHE[5][5] , \CACHE[5][4] ,
         \CACHE[5][3] , \CACHE[5][2] , \CACHE[5][1] , \CACHE[5][0] ,
         \CACHE[4][153] , \CACHE[4][149] , \CACHE[4][148] , \CACHE[4][143] ,
         \CACHE[4][142] , \CACHE[4][141] , \CACHE[4][139] , \CACHE[4][138] ,
         \CACHE[4][137] , \CACHE[4][136] , \CACHE[4][132] , \CACHE[4][131] ,
         \CACHE[4][129] , \CACHE[4][128] , \CACHE[4][127] , \CACHE[4][126] ,
         \CACHE[4][125] , \CACHE[4][124] , \CACHE[4][123] , \CACHE[4][122] ,
         \CACHE[4][121] , \CACHE[4][120] , \CACHE[4][119] , \CACHE[4][118] ,
         \CACHE[4][117] , \CACHE[4][116] , \CACHE[4][115] , \CACHE[4][114] ,
         \CACHE[4][113] , \CACHE[4][112] , \CACHE[4][111] , \CACHE[4][110] ,
         \CACHE[4][109] , \CACHE[4][108] , \CACHE[4][107] , \CACHE[4][106] ,
         \CACHE[4][105] , \CACHE[4][104] , \CACHE[4][103] , \CACHE[4][102] ,
         \CACHE[4][101] , \CACHE[4][100] , \CACHE[4][99] , \CACHE[4][98] ,
         \CACHE[4][97] , \CACHE[4][96] , \CACHE[4][95] , \CACHE[4][94] ,
         \CACHE[4][93] , \CACHE[4][92] , \CACHE[4][91] , \CACHE[4][90] ,
         \CACHE[4][89] , \CACHE[4][88] , \CACHE[4][87] , \CACHE[4][86] ,
         \CACHE[4][85] , \CACHE[4][84] , \CACHE[4][83] , \CACHE[4][82] ,
         \CACHE[4][81] , \CACHE[4][80] , \CACHE[4][79] , \CACHE[4][78] ,
         \CACHE[4][77] , \CACHE[4][76] , \CACHE[4][75] , \CACHE[4][74] ,
         \CACHE[4][73] , \CACHE[4][72] , \CACHE[4][71] , \CACHE[4][70] ,
         \CACHE[4][69] , \CACHE[4][68] , \CACHE[4][67] , \CACHE[4][66] ,
         \CACHE[4][65] , \CACHE[4][64] , \CACHE[4][63] , \CACHE[4][62] ,
         \CACHE[4][61] , \CACHE[4][60] , \CACHE[4][59] , \CACHE[4][58] ,
         \CACHE[4][57] , \CACHE[4][56] , \CACHE[4][55] , \CACHE[4][54] ,
         \CACHE[4][53] , \CACHE[4][52] , \CACHE[4][51] , \CACHE[4][50] ,
         \CACHE[4][49] , \CACHE[4][48] , \CACHE[4][47] , \CACHE[4][46] ,
         \CACHE[4][45] , \CACHE[4][44] , \CACHE[4][43] , \CACHE[4][42] ,
         \CACHE[4][41] , \CACHE[4][40] , \CACHE[4][39] , \CACHE[4][38] ,
         \CACHE[4][37] , \CACHE[4][36] , \CACHE[4][35] , \CACHE[4][34] ,
         \CACHE[4][33] , \CACHE[4][32] , \CACHE[4][31] , \CACHE[4][30] ,
         \CACHE[4][29] , \CACHE[4][28] , \CACHE[4][27] , \CACHE[4][26] ,
         \CACHE[4][25] , \CACHE[4][24] , \CACHE[4][23] , \CACHE[4][22] ,
         \CACHE[4][21] , \CACHE[4][20] , \CACHE[4][19] , \CACHE[4][18] ,
         \CACHE[4][17] , \CACHE[4][16] , \CACHE[4][15] , \CACHE[4][14] ,
         \CACHE[4][13] , \CACHE[4][12] , \CACHE[4][11] , \CACHE[4][10] ,
         \CACHE[4][9] , \CACHE[4][8] , \CACHE[4][7] , \CACHE[4][6] ,
         \CACHE[4][5] , \CACHE[4][4] , \CACHE[4][3] , \CACHE[4][2] ,
         \CACHE[4][1] , \CACHE[4][0] , \CACHE[3][153] , \CACHE[3][149] ,
         \CACHE[3][148] , \CACHE[3][143] , \CACHE[3][142] , \CACHE[3][141] ,
         \CACHE[3][139] , \CACHE[3][138] , \CACHE[3][137] , \CACHE[3][136] ,
         \CACHE[3][135] , \CACHE[3][132] , \CACHE[3][131] , \CACHE[3][129] ,
         \CACHE[3][128] , \CACHE[3][127] , \CACHE[3][126] , \CACHE[3][125] ,
         \CACHE[3][124] , \CACHE[3][123] , \CACHE[3][122] , \CACHE[3][121] ,
         \CACHE[3][120] , \CACHE[3][119] , \CACHE[3][118] , \CACHE[3][117] ,
         \CACHE[3][116] , \CACHE[3][115] , \CACHE[3][114] , \CACHE[3][113] ,
         \CACHE[3][112] , \CACHE[3][111] , \CACHE[3][110] , \CACHE[3][109] ,
         \CACHE[3][108] , \CACHE[3][107] , \CACHE[3][106] , \CACHE[3][105] ,
         \CACHE[3][104] , \CACHE[3][103] , \CACHE[3][102] , \CACHE[3][101] ,
         \CACHE[3][100] , \CACHE[3][99] , \CACHE[3][98] , \CACHE[3][97] ,
         \CACHE[3][96] , \CACHE[3][95] , \CACHE[3][94] , \CACHE[3][93] ,
         \CACHE[3][92] , \CACHE[3][91] , \CACHE[3][90] , \CACHE[3][89] ,
         \CACHE[3][88] , \CACHE[3][87] , \CACHE[3][86] , \CACHE[3][85] ,
         \CACHE[3][84] , \CACHE[3][83] , \CACHE[3][82] , \CACHE[3][81] ,
         \CACHE[3][80] , \CACHE[3][79] , \CACHE[3][78] , \CACHE[3][77] ,
         \CACHE[3][76] , \CACHE[3][75] , \CACHE[3][74] , \CACHE[3][73] ,
         \CACHE[3][72] , \CACHE[3][71] , \CACHE[3][70] , \CACHE[3][69] ,
         \CACHE[3][68] , \CACHE[3][67] , \CACHE[3][66] , \CACHE[3][65] ,
         \CACHE[3][64] , \CACHE[3][63] , \CACHE[3][62] , \CACHE[3][61] ,
         \CACHE[3][60] , \CACHE[3][59] , \CACHE[3][58] , \CACHE[3][57] ,
         \CACHE[3][56] , \CACHE[3][55] , \CACHE[3][54] , \CACHE[3][53] ,
         \CACHE[3][52] , \CACHE[3][51] , \CACHE[3][50] , \CACHE[3][49] ,
         \CACHE[3][48] , \CACHE[3][47] , \CACHE[3][46] , \CACHE[3][45] ,
         \CACHE[3][44] , \CACHE[3][43] , \CACHE[3][42] , \CACHE[3][41] ,
         \CACHE[3][40] , \CACHE[3][39] , \CACHE[3][38] , \CACHE[3][37] ,
         \CACHE[3][36] , \CACHE[3][35] , \CACHE[3][34] , \CACHE[3][33] ,
         \CACHE[3][32] , \CACHE[3][31] , \CACHE[3][30] , \CACHE[3][29] ,
         \CACHE[3][28] , \CACHE[3][27] , \CACHE[3][26] , \CACHE[3][25] ,
         \CACHE[3][24] , \CACHE[3][23] , \CACHE[3][22] , \CACHE[3][21] ,
         \CACHE[3][20] , \CACHE[3][19] , \CACHE[3][18] , \CACHE[3][17] ,
         \CACHE[3][16] , \CACHE[3][15] , \CACHE[3][14] , \CACHE[3][13] ,
         \CACHE[3][12] , \CACHE[3][11] , \CACHE[3][10] , \CACHE[3][9] ,
         \CACHE[3][8] , \CACHE[3][7] , \CACHE[3][6] , \CACHE[3][5] ,
         \CACHE[3][4] , \CACHE[3][3] , \CACHE[3][2] , \CACHE[3][1] ,
         \CACHE[3][0] , \CACHE[2][153] , \CACHE[2][149] , \CACHE[2][148] ,
         \CACHE[2][143] , \CACHE[2][142] , \CACHE[2][141] , \CACHE[2][139] ,
         \CACHE[2][138] , \CACHE[2][137] , \CACHE[2][136] , \CACHE[2][135] ,
         \CACHE[2][132] , \CACHE[2][131] , \CACHE[2][129] , \CACHE[2][128] ,
         \CACHE[2][127] , \CACHE[2][126] , \CACHE[2][125] , \CACHE[2][124] ,
         \CACHE[2][123] , \CACHE[2][122] , \CACHE[2][121] , \CACHE[2][120] ,
         \CACHE[2][119] , \CACHE[2][118] , \CACHE[2][117] , \CACHE[2][116] ,
         \CACHE[2][115] , \CACHE[2][114] , \CACHE[2][113] , \CACHE[2][112] ,
         \CACHE[2][111] , \CACHE[2][110] , \CACHE[2][109] , \CACHE[2][108] ,
         \CACHE[2][107] , \CACHE[2][106] , \CACHE[2][105] , \CACHE[2][104] ,
         \CACHE[2][103] , \CACHE[2][102] , \CACHE[2][101] , \CACHE[2][100] ,
         \CACHE[2][99] , \CACHE[2][98] , \CACHE[2][97] , \CACHE[2][96] ,
         \CACHE[2][95] , \CACHE[2][94] , \CACHE[2][93] , \CACHE[2][92] ,
         \CACHE[2][91] , \CACHE[2][90] , \CACHE[2][89] , \CACHE[2][88] ,
         \CACHE[2][87] , \CACHE[2][86] , \CACHE[2][85] , \CACHE[2][84] ,
         \CACHE[2][83] , \CACHE[2][82] , \CACHE[2][81] , \CACHE[2][80] ,
         \CACHE[2][79] , \CACHE[2][78] , \CACHE[2][77] , \CACHE[2][76] ,
         \CACHE[2][75] , \CACHE[2][74] , \CACHE[2][73] , \CACHE[2][72] ,
         \CACHE[2][71] , \CACHE[2][70] , \CACHE[2][69] , \CACHE[2][68] ,
         \CACHE[2][67] , \CACHE[2][66] , \CACHE[2][65] , \CACHE[2][64] ,
         \CACHE[2][63] , \CACHE[2][62] , \CACHE[2][61] , \CACHE[2][60] ,
         \CACHE[2][59] , \CACHE[2][58] , \CACHE[2][57] , \CACHE[2][56] ,
         \CACHE[2][55] , \CACHE[2][54] , \CACHE[2][53] , \CACHE[2][52] ,
         \CACHE[2][51] , \CACHE[2][50] , \CACHE[2][49] , \CACHE[2][48] ,
         \CACHE[2][47] , \CACHE[2][46] , \CACHE[2][45] , \CACHE[2][44] ,
         \CACHE[2][43] , \CACHE[2][42] , \CACHE[2][41] , \CACHE[2][40] ,
         \CACHE[2][39] , \CACHE[2][38] , \CACHE[2][37] , \CACHE[2][36] ,
         \CACHE[2][35] , \CACHE[2][34] , \CACHE[2][33] , \CACHE[2][32] ,
         \CACHE[2][31] , \CACHE[2][30] , \CACHE[2][29] , \CACHE[2][28] ,
         \CACHE[2][27] , \CACHE[2][26] , \CACHE[2][25] , \CACHE[2][24] ,
         \CACHE[2][23] , \CACHE[2][22] , \CACHE[2][21] , \CACHE[2][20] ,
         \CACHE[2][19] , \CACHE[2][18] , \CACHE[2][17] , \CACHE[2][16] ,
         \CACHE[2][15] , \CACHE[2][14] , \CACHE[2][13] , \CACHE[2][12] ,
         \CACHE[2][11] , \CACHE[2][10] , \CACHE[2][9] , \CACHE[2][8] ,
         \CACHE[2][7] , \CACHE[2][6] , \CACHE[2][5] , \CACHE[2][4] ,
         \CACHE[2][3] , \CACHE[2][2] , \CACHE[2][1] , \CACHE[2][0] ,
         \CACHE[1][153] , \CACHE[1][149] , \CACHE[1][148] , \CACHE[1][143] ,
         \CACHE[1][142] , \CACHE[1][141] , \CACHE[1][139] , \CACHE[1][138] ,
         \CACHE[1][137] , \CACHE[1][136] , \CACHE[1][135] , \CACHE[1][132] ,
         \CACHE[1][131] , \CACHE[1][129] , \CACHE[1][128] , \CACHE[1][127] ,
         \CACHE[1][126] , \CACHE[1][125] , \CACHE[1][124] , \CACHE[1][123] ,
         \CACHE[1][122] , \CACHE[1][121] , \CACHE[1][120] , \CACHE[1][119] ,
         \CACHE[1][118] , \CACHE[1][117] , \CACHE[1][116] , \CACHE[1][115] ,
         \CACHE[1][114] , \CACHE[1][113] , \CACHE[1][112] , \CACHE[1][111] ,
         \CACHE[1][110] , \CACHE[1][109] , \CACHE[1][108] , \CACHE[1][107] ,
         \CACHE[1][106] , \CACHE[1][105] , \CACHE[1][104] , \CACHE[1][103] ,
         \CACHE[1][102] , \CACHE[1][101] , \CACHE[1][100] , \CACHE[1][99] ,
         \CACHE[1][98] , \CACHE[1][97] , \CACHE[1][96] , \CACHE[1][95] ,
         \CACHE[1][94] , \CACHE[1][93] , \CACHE[1][92] , \CACHE[1][91] ,
         \CACHE[1][90] , \CACHE[1][89] , \CACHE[1][88] , \CACHE[1][87] ,
         \CACHE[1][86] , \CACHE[1][85] , \CACHE[1][84] , \CACHE[1][83] ,
         \CACHE[1][82] , \CACHE[1][81] , \CACHE[1][80] , \CACHE[1][79] ,
         \CACHE[1][78] , \CACHE[1][77] , \CACHE[1][76] , \CACHE[1][75] ,
         \CACHE[1][74] , \CACHE[1][73] , \CACHE[1][72] , \CACHE[1][71] ,
         \CACHE[1][70] , \CACHE[1][69] , \CACHE[1][68] , \CACHE[1][67] ,
         \CACHE[1][66] , \CACHE[1][65] , \CACHE[1][64] , \CACHE[1][63] ,
         \CACHE[1][62] , \CACHE[1][61] , \CACHE[1][60] , \CACHE[1][59] ,
         \CACHE[1][58] , \CACHE[1][57] , \CACHE[1][56] , \CACHE[1][55] ,
         \CACHE[1][54] , \CACHE[1][53] , \CACHE[1][52] , \CACHE[1][51] ,
         \CACHE[1][50] , \CACHE[1][49] , \CACHE[1][48] , \CACHE[1][47] ,
         \CACHE[1][46] , \CACHE[1][45] , \CACHE[1][44] , \CACHE[1][43] ,
         \CACHE[1][42] , \CACHE[1][41] , \CACHE[1][40] , \CACHE[1][39] ,
         \CACHE[1][38] , \CACHE[1][37] , \CACHE[1][36] , \CACHE[1][35] ,
         \CACHE[1][34] , \CACHE[1][33] , \CACHE[1][32] , \CACHE[1][31] ,
         \CACHE[1][30] , \CACHE[1][29] , \CACHE[1][28] , \CACHE[1][27] ,
         \CACHE[1][26] , \CACHE[1][25] , \CACHE[1][24] , \CACHE[1][23] ,
         \CACHE[1][22] , \CACHE[1][21] , \CACHE[1][20] , \CACHE[1][19] ,
         \CACHE[1][18] , \CACHE[1][17] , \CACHE[1][16] , \CACHE[1][15] ,
         \CACHE[1][14] , \CACHE[1][13] , \CACHE[1][12] , \CACHE[1][11] ,
         \CACHE[1][10] , \CACHE[1][9] , \CACHE[1][8] , \CACHE[1][7] ,
         \CACHE[1][6] , \CACHE[1][5] , \CACHE[1][4] , \CACHE[1][3] ,
         \CACHE[1][2] , \CACHE[1][1] , \CACHE[1][0] , \CACHE[0][153] ,
         \CACHE[0][149] , \CACHE[0][148] , \CACHE[0][143] , \CACHE[0][142] ,
         \CACHE[0][141] , \CACHE[0][139] , \CACHE[0][138] , \CACHE[0][137] ,
         \CACHE[0][136] , \CACHE[0][135] , \CACHE[0][132] , \CACHE[0][131] ,
         \CACHE[0][129] , \CACHE[0][128] , \CACHE[0][127] , \CACHE[0][126] ,
         \CACHE[0][125] , \CACHE[0][124] , \CACHE[0][123] , \CACHE[0][122] ,
         \CACHE[0][121] , \CACHE[0][120] , \CACHE[0][119] , \CACHE[0][118] ,
         \CACHE[0][117] , \CACHE[0][116] , \CACHE[0][115] , \CACHE[0][114] ,
         \CACHE[0][113] , \CACHE[0][112] , \CACHE[0][111] , \CACHE[0][110] ,
         \CACHE[0][109] , \CACHE[0][108] , \CACHE[0][107] , \CACHE[0][106] ,
         \CACHE[0][105] , \CACHE[0][104] , \CACHE[0][103] , \CACHE[0][102] ,
         \CACHE[0][101] , \CACHE[0][100] , \CACHE[0][99] , \CACHE[0][98] ,
         \CACHE[0][97] , \CACHE[0][96] , \CACHE[0][95] , \CACHE[0][94] ,
         \CACHE[0][93] , \CACHE[0][92] , \CACHE[0][91] , \CACHE[0][90] ,
         \CACHE[0][89] , \CACHE[0][88] , \CACHE[0][87] , \CACHE[0][86] ,
         \CACHE[0][85] , \CACHE[0][84] , \CACHE[0][83] , \CACHE[0][82] ,
         \CACHE[0][81] , \CACHE[0][80] , \CACHE[0][79] , \CACHE[0][78] ,
         \CACHE[0][77] , \CACHE[0][76] , \CACHE[0][75] , \CACHE[0][74] ,
         \CACHE[0][73] , \CACHE[0][72] , \CACHE[0][71] , \CACHE[0][70] ,
         \CACHE[0][69] , \CACHE[0][68] , \CACHE[0][67] , \CACHE[0][66] ,
         \CACHE[0][65] , \CACHE[0][64] , \CACHE[0][63] , \CACHE[0][62] ,
         \CACHE[0][61] , \CACHE[0][60] , \CACHE[0][59] , \CACHE[0][58] ,
         \CACHE[0][57] , \CACHE[0][56] , \CACHE[0][55] , \CACHE[0][54] ,
         \CACHE[0][53] , \CACHE[0][52] , \CACHE[0][51] , \CACHE[0][50] ,
         \CACHE[0][49] , \CACHE[0][48] , \CACHE[0][47] , \CACHE[0][46] ,
         \CACHE[0][45] , \CACHE[0][44] , \CACHE[0][43] , \CACHE[0][42] ,
         \CACHE[0][41] , \CACHE[0][40] , \CACHE[0][39] , \CACHE[0][38] ,
         \CACHE[0][37] , \CACHE[0][36] , \CACHE[0][35] , \CACHE[0][34] ,
         \CACHE[0][33] , \CACHE[0][32] , \CACHE[0][31] , \CACHE[0][30] ,
         \CACHE[0][29] , \CACHE[0][28] , \CACHE[0][27] , \CACHE[0][26] ,
         \CACHE[0][25] , \CACHE[0][24] , \CACHE[0][23] , \CACHE[0][22] ,
         \CACHE[0][21] , \CACHE[0][20] , \CACHE[0][19] , \CACHE[0][18] ,
         \CACHE[0][17] , \CACHE[0][16] , \CACHE[0][15] , \CACHE[0][14] ,
         \CACHE[0][13] , \CACHE[0][12] , \CACHE[0][11] , \CACHE[0][10] ,
         \CACHE[0][9] , \CACHE[0][8] , \CACHE[0][7] , \CACHE[0][6] ,
         \CACHE[0][5] , \CACHE[0][4] , \CACHE[0][3] , \CACHE[0][2] ,
         \CACHE[0][1] , \CACHE[0][0] , N33, N34, N35, N36, N37, N38, N40, N41,
         N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, n7, n8, n10, n12, n14, n15, n17, n21, n26, n31,
         n36, n41, n46, n51, n56, n61, n66, n71, n76, n81, n86, n91, n96, n101,
         n106, n111, n116, n121, n126, n131, n136, n141, n146, n151, n156,
         n161, n166, n171, n176, n177, n178, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n338, n341, n343, n345,
         n347, n349, n351, n352, n353, n355, n356, n358, n359, n361, n362,
         n363, n364, n365, n366, n368, n369, n371, n373, n375, n377, n379,
         n381, n383, n385, n387, n389, n395, n397, n399, n401, n403, n407,
         n409, n411, n413, n415, n417, n419, n421, n423, n425, n427, n428,
         n429, n430, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178;
  assign N30 = proc_addr[2];
  assign N31 = proc_addr[3];
  assign N32 = proc_addr[4];

  DFFRX1 \CACHE_reg[7][118]  ( .D(n3015), .CK(clk), .RN(n3834), .Q(
        \CACHE[7][118] ), .QN(n1775) );
  DFFRX1 \CACHE_reg[7][117]  ( .D(n3014), .CK(clk), .RN(n3834), .Q(
        \CACHE[7][117] ), .QN(n1774) );
  DFFRX1 \CACHE_reg[7][116]  ( .D(n3013), .CK(clk), .RN(n3834), .Q(
        \CACHE[7][116] ), .QN(n1773) );
  DFFRX1 \CACHE_reg[7][115]  ( .D(n3012), .CK(clk), .RN(n3834), .Q(
        \CACHE[7][115] ), .QN(n1772) );
  DFFRX1 \CACHE_reg[7][114]  ( .D(n3011), .CK(clk), .RN(n3833), .Q(
        \CACHE[7][114] ), .QN(n1771) );
  DFFRX1 \CACHE_reg[7][113]  ( .D(n3010), .CK(clk), .RN(n3833), .Q(
        \CACHE[7][113] ), .QN(n1770) );
  DFFRX1 \CACHE_reg[7][112]  ( .D(n3009), .CK(clk), .RN(n3833), .Q(
        \CACHE[7][112] ), .QN(n1769) );
  DFFRX1 \CACHE_reg[7][111]  ( .D(n3008), .CK(clk), .RN(n3833), .Q(
        \CACHE[7][111] ), .QN(n1768) );
  DFFRX1 \CACHE_reg[7][110]  ( .D(n3007), .CK(clk), .RN(n3833), .Q(
        \CACHE[7][110] ), .QN(n1767) );
  DFFRX1 \CACHE_reg[7][109]  ( .D(n3006), .CK(clk), .RN(n3833), .Q(
        \CACHE[7][109] ), .QN(n1766) );
  DFFRX1 \CACHE_reg[7][108]  ( .D(n3005), .CK(clk), .RN(n3833), .Q(
        \CACHE[7][108] ), .QN(n1765) );
  DFFRX1 \CACHE_reg[7][107]  ( .D(n3004), .CK(clk), .RN(n3833), .Q(
        \CACHE[7][107] ), .QN(n1764) );
  DFFRX1 \CACHE_reg[7][106]  ( .D(n3003), .CK(clk), .RN(n3833), .Q(
        \CACHE[7][106] ), .QN(n1763) );
  DFFRX1 \CACHE_reg[7][105]  ( .D(n3002), .CK(clk), .RN(n3833), .Q(
        \CACHE[7][105] ), .QN(n1762) );
  DFFRX1 \CACHE_reg[7][104]  ( .D(n3001), .CK(clk), .RN(n3833), .Q(
        \CACHE[7][104] ), .QN(n1761) );
  DFFRX1 \CACHE_reg[7][103]  ( .D(n3000), .CK(clk), .RN(n3833), .Q(
        \CACHE[7][103] ), .QN(n1760) );
  DFFRX1 \CACHE_reg[7][102]  ( .D(n2999), .CK(clk), .RN(n3832), .Q(
        \CACHE[7][102] ), .QN(n1759) );
  DFFRX1 \CACHE_reg[7][101]  ( .D(n2998), .CK(clk), .RN(n3832), .Q(
        \CACHE[7][101] ), .QN(n1758) );
  DFFRX1 \CACHE_reg[7][100]  ( .D(n2997), .CK(clk), .RN(n3832), .Q(
        \CACHE[7][100] ), .QN(n1757) );
  DFFRX1 \CACHE_reg[7][99]  ( .D(n2996), .CK(clk), .RN(n3832), .Q(
        \CACHE[7][99] ), .QN(n1756) );
  DFFRX1 \CACHE_reg[7][98]  ( .D(n2995), .CK(clk), .RN(n3832), .Q(
        \CACHE[7][98] ), .QN(n1755) );
  DFFRX1 \CACHE_reg[7][97]  ( .D(n2994), .CK(clk), .RN(n3832), .Q(
        \CACHE[7][97] ), .QN(n1754) );
  DFFRX1 \CACHE_reg[7][96]  ( .D(n2993), .CK(clk), .RN(n3832), .Q(
        \CACHE[7][96] ), .QN(n1753) );
  DFFRX1 \CACHE_reg[7][95]  ( .D(n2992), .CK(clk), .RN(n3832), .Q(
        \CACHE[7][95] ), .QN(n1752) );
  DFFRX1 \CACHE_reg[7][94]  ( .D(n2991), .CK(clk), .RN(n3832), .Q(
        \CACHE[7][94] ), .QN(n1751) );
  DFFRX1 \CACHE_reg[7][93]  ( .D(n2990), .CK(clk), .RN(n3832), .Q(
        \CACHE[7][93] ), .QN(n1750) );
  DFFRX1 \CACHE_reg[7][92]  ( .D(n2989), .CK(clk), .RN(n3832), .Q(
        \CACHE[7][92] ), .QN(n1749) );
  DFFRX1 \CACHE_reg[7][91]  ( .D(n2988), .CK(clk), .RN(n3832), .Q(
        \CACHE[7][91] ), .QN(n1748) );
  DFFRX1 \CACHE_reg[7][90]  ( .D(n2987), .CK(clk), .RN(n3831), .Q(
        \CACHE[7][90] ), .QN(n1747) );
  DFFRX1 \CACHE_reg[7][89]  ( .D(n2986), .CK(clk), .RN(n3831), .Q(
        \CACHE[7][89] ), .QN(n1746) );
  DFFRX1 \CACHE_reg[7][88]  ( .D(n2985), .CK(clk), .RN(n3831), .Q(
        \CACHE[7][88] ), .QN(n1745) );
  DFFRX1 \CACHE_reg[7][87]  ( .D(n2984), .CK(clk), .RN(n3831), .Q(
        \CACHE[7][87] ), .QN(n1744) );
  DFFRX1 \CACHE_reg[7][86]  ( .D(n2983), .CK(clk), .RN(n3831), .Q(
        \CACHE[7][86] ), .QN(n1743) );
  DFFRX1 \CACHE_reg[7][85]  ( .D(n2982), .CK(clk), .RN(n3831), .Q(
        \CACHE[7][85] ), .QN(n1742) );
  DFFRX1 \CACHE_reg[7][84]  ( .D(n2981), .CK(clk), .RN(n3831), .Q(
        \CACHE[7][84] ), .QN(n1741) );
  DFFRX1 \CACHE_reg[7][83]  ( .D(n2980), .CK(clk), .RN(n3831), .Q(
        \CACHE[7][83] ), .QN(n1740) );
  DFFRX1 \CACHE_reg[7][82]  ( .D(n2979), .CK(clk), .RN(n3831), .Q(
        \CACHE[7][82] ), .QN(n1739) );
  DFFRX1 \CACHE_reg[7][81]  ( .D(n2978), .CK(clk), .RN(n3831), .Q(
        \CACHE[7][81] ), .QN(n1738) );
  DFFRX1 \CACHE_reg[7][80]  ( .D(n2977), .CK(clk), .RN(n3831), .Q(
        \CACHE[7][80] ), .QN(n1737) );
  DFFRX1 \CACHE_reg[7][79]  ( .D(n2976), .CK(clk), .RN(n3831), .Q(
        \CACHE[7][79] ), .QN(n1736) );
  DFFRX1 \CACHE_reg[7][78]  ( .D(n2975), .CK(clk), .RN(n3830), .Q(
        \CACHE[7][78] ), .QN(n1735) );
  DFFRX1 \CACHE_reg[7][77]  ( .D(n2974), .CK(clk), .RN(n3830), .Q(
        \CACHE[7][77] ), .QN(n1734) );
  DFFRX1 \CACHE_reg[7][76]  ( .D(n2973), .CK(clk), .RN(n3830), .Q(
        \CACHE[7][76] ), .QN(n1733) );
  DFFRX1 \CACHE_reg[7][75]  ( .D(n2972), .CK(clk), .RN(n3830), .Q(
        \CACHE[7][75] ), .QN(n1732) );
  DFFRX1 \CACHE_reg[7][74]  ( .D(n2971), .CK(clk), .RN(n3830), .Q(
        \CACHE[7][74] ), .QN(n1731) );
  DFFRX1 \CACHE_reg[7][73]  ( .D(n2970), .CK(clk), .RN(n3830), .Q(
        \CACHE[7][73] ), .QN(n1730) );
  DFFRX1 \CACHE_reg[7][72]  ( .D(n2969), .CK(clk), .RN(n3830), .Q(
        \CACHE[7][72] ), .QN(n1729) );
  DFFRX1 \CACHE_reg[7][71]  ( .D(n2968), .CK(clk), .RN(n3830), .Q(
        \CACHE[7][71] ), .QN(n1728) );
  DFFRX1 \CACHE_reg[7][70]  ( .D(n2967), .CK(clk), .RN(n3830), .Q(
        \CACHE[7][70] ), .QN(n1727) );
  DFFRX1 \CACHE_reg[7][69]  ( .D(n2966), .CK(clk), .RN(n3830), .Q(
        \CACHE[7][69] ), .QN(n1726) );
  DFFRX1 \CACHE_reg[7][68]  ( .D(n2965), .CK(clk), .RN(n3830), .Q(
        \CACHE[7][68] ), .QN(n1725) );
  DFFRX1 \CACHE_reg[7][67]  ( .D(n2964), .CK(clk), .RN(n3830), .Q(
        \CACHE[7][67] ), .QN(n1724) );
  DFFRX1 \CACHE_reg[7][66]  ( .D(n2963), .CK(clk), .RN(n3829), .Q(
        \CACHE[7][66] ), .QN(n1723) );
  DFFRX1 \CACHE_reg[7][65]  ( .D(n2962), .CK(clk), .RN(n3829), .Q(
        \CACHE[7][65] ), .QN(n1722) );
  DFFRX1 \CACHE_reg[7][64]  ( .D(n2961), .CK(clk), .RN(n3829), .Q(
        \CACHE[7][64] ), .QN(n1721) );
  DFFRX1 \CACHE_reg[7][63]  ( .D(n2960), .CK(clk), .RN(n3829), .Q(
        \CACHE[7][63] ), .QN(n1720) );
  DFFRX1 \CACHE_reg[7][62]  ( .D(n2959), .CK(clk), .RN(n3829), .Q(
        \CACHE[7][62] ), .QN(n1719) );
  DFFRX1 \CACHE_reg[7][61]  ( .D(n2958), .CK(clk), .RN(n3829), .Q(
        \CACHE[7][61] ), .QN(n1718) );
  DFFRX1 \CACHE_reg[7][60]  ( .D(n2957), .CK(clk), .RN(n3829), .Q(
        \CACHE[7][60] ), .QN(n1717) );
  DFFRX1 \CACHE_reg[7][59]  ( .D(n2956), .CK(clk), .RN(n3829), .Q(
        \CACHE[7][59] ), .QN(n1716) );
  DFFRX1 \CACHE_reg[7][58]  ( .D(n2955), .CK(clk), .RN(n3829), .Q(
        \CACHE[7][58] ), .QN(n1715) );
  DFFRX1 \CACHE_reg[7][57]  ( .D(n2954), .CK(clk), .RN(n3829), .Q(
        \CACHE[7][57] ), .QN(n1714) );
  DFFRX1 \CACHE_reg[7][56]  ( .D(n2953), .CK(clk), .RN(n3829), .Q(
        \CACHE[7][56] ), .QN(n1713) );
  DFFRX1 \CACHE_reg[7][55]  ( .D(n2952), .CK(clk), .RN(n3829), .Q(
        \CACHE[7][55] ), .QN(n1712) );
  DFFRX1 \CACHE_reg[7][54]  ( .D(n2951), .CK(clk), .RN(n3828), .Q(
        \CACHE[7][54] ), .QN(n1711) );
  DFFRX1 \CACHE_reg[7][53]  ( .D(n2950), .CK(clk), .RN(n3828), .Q(
        \CACHE[7][53] ), .QN(n1710) );
  DFFRX1 \CACHE_reg[7][52]  ( .D(n2949), .CK(clk), .RN(n3828), .Q(
        \CACHE[7][52] ), .QN(n1709) );
  DFFRX1 \CACHE_reg[7][51]  ( .D(n2948), .CK(clk), .RN(n3828), .Q(
        \CACHE[7][51] ), .QN(n1708) );
  DFFRX1 \CACHE_reg[7][50]  ( .D(n2947), .CK(clk), .RN(n3828), .Q(
        \CACHE[7][50] ), .QN(n1707) );
  DFFRX1 \CACHE_reg[7][49]  ( .D(n2946), .CK(clk), .RN(n3828), .Q(
        \CACHE[7][49] ), .QN(n1706) );
  DFFRX1 \CACHE_reg[7][48]  ( .D(n2945), .CK(clk), .RN(n3828), .Q(
        \CACHE[7][48] ), .QN(n1705) );
  DFFRX1 \CACHE_reg[7][47]  ( .D(n2944), .CK(clk), .RN(n3828), .Q(
        \CACHE[7][47] ), .QN(n1704) );
  DFFRX1 \CACHE_reg[7][46]  ( .D(n2943), .CK(clk), .RN(n3828), .Q(
        \CACHE[7][46] ), .QN(n1703) );
  DFFRX1 \CACHE_reg[7][45]  ( .D(n2942), .CK(clk), .RN(n3828), .Q(
        \CACHE[7][45] ), .QN(n1702) );
  DFFRX1 \CACHE_reg[7][44]  ( .D(n2941), .CK(clk), .RN(n3828), .Q(
        \CACHE[7][44] ), .QN(n1701) );
  DFFRX1 \CACHE_reg[7][43]  ( .D(n2940), .CK(clk), .RN(n3828), .Q(
        \CACHE[7][43] ), .QN(n1700) );
  DFFRX1 \CACHE_reg[7][42]  ( .D(n2939), .CK(clk), .RN(n3827), .Q(
        \CACHE[7][42] ), .QN(n1699) );
  DFFRX1 \CACHE_reg[7][41]  ( .D(n2938), .CK(clk), .RN(n3827), .Q(
        \CACHE[7][41] ), .QN(n1698) );
  DFFRX1 \CACHE_reg[7][40]  ( .D(n2937), .CK(clk), .RN(n3827), .Q(
        \CACHE[7][40] ), .QN(n1697) );
  DFFRX1 \CACHE_reg[7][39]  ( .D(n2936), .CK(clk), .RN(n3827), .Q(
        \CACHE[7][39] ), .QN(n1696) );
  DFFRX1 \CACHE_reg[7][38]  ( .D(n2935), .CK(clk), .RN(n3827), .Q(
        \CACHE[7][38] ), .QN(n1695) );
  DFFRX1 \CACHE_reg[7][37]  ( .D(n2934), .CK(clk), .RN(n3827), .Q(
        \CACHE[7][37] ), .QN(n1694) );
  DFFRX1 \CACHE_reg[7][36]  ( .D(n2933), .CK(clk), .RN(n3827), .Q(
        \CACHE[7][36] ), .QN(n1693) );
  DFFRX1 \CACHE_reg[7][35]  ( .D(n2932), .CK(clk), .RN(n3827), .Q(
        \CACHE[7][35] ), .QN(n1692) );
  DFFRX1 \CACHE_reg[7][34]  ( .D(n2931), .CK(clk), .RN(n3827), .Q(
        \CACHE[7][34] ), .QN(n1691) );
  DFFRX1 \CACHE_reg[7][33]  ( .D(n2930), .CK(clk), .RN(n3827), .Q(
        \CACHE[7][33] ), .QN(n1690) );
  DFFRX1 \CACHE_reg[7][32]  ( .D(n2929), .CK(clk), .RN(n3827), .Q(
        \CACHE[7][32] ), .QN(n1689) );
  DFFRX1 \CACHE_reg[7][31]  ( .D(n2928), .CK(clk), .RN(n3827), .Q(
        \CACHE[7][31] ), .QN(n1688) );
  DFFRX1 \CACHE_reg[7][30]  ( .D(n2927), .CK(clk), .RN(n3826), .Q(
        \CACHE[7][30] ), .QN(n1687) );
  DFFRX1 \CACHE_reg[7][29]  ( .D(n2926), .CK(clk), .RN(n3826), .Q(
        \CACHE[7][29] ), .QN(n1686) );
  DFFRX1 \CACHE_reg[7][28]  ( .D(n2925), .CK(clk), .RN(n3826), .Q(
        \CACHE[7][28] ), .QN(n1685) );
  DFFRX1 \CACHE_reg[7][27]  ( .D(n2924), .CK(clk), .RN(n3826), .Q(
        \CACHE[7][27] ), .QN(n1684) );
  DFFRX1 \CACHE_reg[7][26]  ( .D(n2923), .CK(clk), .RN(n3826), .Q(
        \CACHE[7][26] ), .QN(n1683) );
  DFFRX1 \CACHE_reg[7][25]  ( .D(n2922), .CK(clk), .RN(n3826), .Q(
        \CACHE[7][25] ), .QN(n1682) );
  DFFRX1 \CACHE_reg[7][24]  ( .D(n2921), .CK(clk), .RN(n3826), .Q(
        \CACHE[7][24] ), .QN(n1681) );
  DFFRX1 \CACHE_reg[7][23]  ( .D(n2920), .CK(clk), .RN(n3826), .Q(
        \CACHE[7][23] ), .QN(n1680) );
  DFFRX1 \CACHE_reg[7][22]  ( .D(n2919), .CK(clk), .RN(n3826), .Q(
        \CACHE[7][22] ), .QN(n1679) );
  DFFRX1 \CACHE_reg[7][21]  ( .D(n2918), .CK(clk), .RN(n3826), .Q(
        \CACHE[7][21] ), .QN(n1678) );
  DFFRX1 \CACHE_reg[7][20]  ( .D(n2917), .CK(clk), .RN(n3826), .Q(
        \CACHE[7][20] ), .QN(n1677) );
  DFFRX1 \CACHE_reg[7][19]  ( .D(n2916), .CK(clk), .RN(n3826), .Q(
        \CACHE[7][19] ), .QN(n1676) );
  DFFRX1 \CACHE_reg[7][18]  ( .D(n2915), .CK(clk), .RN(n3825), .Q(
        \CACHE[7][18] ), .QN(n1675) );
  DFFRX1 \CACHE_reg[7][17]  ( .D(n2914), .CK(clk), .RN(n3825), .Q(
        \CACHE[7][17] ), .QN(n1674) );
  DFFRX1 \CACHE_reg[7][16]  ( .D(n2913), .CK(clk), .RN(n3825), .Q(
        \CACHE[7][16] ), .QN(n1673) );
  DFFRX1 \CACHE_reg[7][15]  ( .D(n2912), .CK(clk), .RN(n3825), .Q(
        \CACHE[7][15] ), .QN(n1672) );
  DFFRX1 \CACHE_reg[7][14]  ( .D(n2911), .CK(clk), .RN(n3825), .Q(
        \CACHE[7][14] ), .QN(n1671) );
  DFFRX1 \CACHE_reg[7][13]  ( .D(n2910), .CK(clk), .RN(n3825), .Q(
        \CACHE[7][13] ), .QN(n1670) );
  DFFRX1 \CACHE_reg[7][12]  ( .D(n2909), .CK(clk), .RN(n3825), .Q(
        \CACHE[7][12] ), .QN(n1669) );
  DFFRX1 \CACHE_reg[7][11]  ( .D(n2908), .CK(clk), .RN(n3825), .Q(
        \CACHE[7][11] ), .QN(n1668) );
  DFFRX1 \CACHE_reg[7][10]  ( .D(n2907), .CK(clk), .RN(n3825), .Q(
        \CACHE[7][10] ), .QN(n1667) );
  DFFRX1 \CACHE_reg[7][9]  ( .D(n2906), .CK(clk), .RN(n3825), .Q(\CACHE[7][9] ), .QN(n1666) );
  DFFRX1 \CACHE_reg[7][8]  ( .D(n2905), .CK(clk), .RN(n3825), .Q(\CACHE[7][8] ), .QN(n1665) );
  DFFRX1 \CACHE_reg[7][7]  ( .D(n2904), .CK(clk), .RN(n3825), .Q(\CACHE[7][7] ), .QN(n1664) );
  DFFRX1 \CACHE_reg[7][6]  ( .D(n2903), .CK(clk), .RN(n3824), .Q(\CACHE[7][6] ), .QN(n1663) );
  DFFRX1 \CACHE_reg[7][5]  ( .D(n2902), .CK(clk), .RN(n3824), .Q(\CACHE[7][5] ), .QN(n1662) );
  DFFRX1 \CACHE_reg[7][4]  ( .D(n2901), .CK(clk), .RN(n3824), .Q(\CACHE[7][4] ), .QN(n1661) );
  DFFRX1 \CACHE_reg[7][3]  ( .D(n2900), .CK(clk), .RN(n3824), .Q(\CACHE[7][3] ), .QN(n1660) );
  DFFRX1 \CACHE_reg[7][2]  ( .D(n2899), .CK(clk), .RN(n3824), .Q(\CACHE[7][2] ), .QN(n1659) );
  DFFRX1 \CACHE_reg[7][1]  ( .D(n2898), .CK(clk), .RN(n3824), .Q(\CACHE[7][1] ), .QN(n1658) );
  DFFRX1 \CACHE_reg[7][0]  ( .D(n2897), .CK(clk), .RN(n3824), .Q(\CACHE[7][0] ), .QN(n1657) );
  DFFRX1 \CACHE_reg[3][118]  ( .D(n2395), .CK(clk), .RN(n3782), .Q(
        \CACHE[3][118] ), .QN(n1155) );
  DFFRX1 \CACHE_reg[3][117]  ( .D(n2394), .CK(clk), .RN(n3782), .Q(
        \CACHE[3][117] ), .QN(n1154) );
  DFFRX1 \CACHE_reg[3][116]  ( .D(n2393), .CK(clk), .RN(n3782), .Q(
        \CACHE[3][116] ), .QN(n1153) );
  DFFRX1 \CACHE_reg[3][115]  ( .D(n2392), .CK(clk), .RN(n3782), .Q(
        \CACHE[3][115] ), .QN(n1152) );
  DFFRX1 \CACHE_reg[3][114]  ( .D(n2391), .CK(clk), .RN(n3782), .Q(
        \CACHE[3][114] ), .QN(n1151) );
  DFFRX1 \CACHE_reg[3][113]  ( .D(n2390), .CK(clk), .RN(n3782), .Q(
        \CACHE[3][113] ), .QN(n1150) );
  DFFRX1 \CACHE_reg[3][112]  ( .D(n2389), .CK(clk), .RN(n3782), .Q(
        \CACHE[3][112] ), .QN(n1149) );
  DFFRX1 \CACHE_reg[3][111]  ( .D(n2388), .CK(clk), .RN(n3782), .Q(
        \CACHE[3][111] ), .QN(n1148) );
  DFFRX1 \CACHE_reg[3][110]  ( .D(n2387), .CK(clk), .RN(n3781), .Q(
        \CACHE[3][110] ), .QN(n1147) );
  DFFRX1 \CACHE_reg[3][109]  ( .D(n2386), .CK(clk), .RN(n3781), .Q(
        \CACHE[3][109] ), .QN(n1146) );
  DFFRX1 \CACHE_reg[3][108]  ( .D(n2385), .CK(clk), .RN(n3781), .Q(
        \CACHE[3][108] ), .QN(n1145) );
  DFFRX1 \CACHE_reg[3][107]  ( .D(n2384), .CK(clk), .RN(n3781), .Q(
        \CACHE[3][107] ), .QN(n1144) );
  DFFRX1 \CACHE_reg[3][106]  ( .D(n2383), .CK(clk), .RN(n3781), .Q(
        \CACHE[3][106] ), .QN(n1143) );
  DFFRX1 \CACHE_reg[3][105]  ( .D(n2382), .CK(clk), .RN(n3781), .Q(
        \CACHE[3][105] ), .QN(n1142) );
  DFFRX1 \CACHE_reg[3][104]  ( .D(n2381), .CK(clk), .RN(n3781), .Q(
        \CACHE[3][104] ), .QN(n1141) );
  DFFRX1 \CACHE_reg[3][103]  ( .D(n2380), .CK(clk), .RN(n3781), .Q(
        \CACHE[3][103] ), .QN(n1140) );
  DFFRX1 \CACHE_reg[3][102]  ( .D(n2379), .CK(clk), .RN(n3781), .Q(
        \CACHE[3][102] ), .QN(n1139) );
  DFFRX1 \CACHE_reg[3][101]  ( .D(n2378), .CK(clk), .RN(n3781), .Q(
        \CACHE[3][101] ), .QN(n1138) );
  DFFRX1 \CACHE_reg[3][100]  ( .D(n2377), .CK(clk), .RN(n3781), .Q(
        \CACHE[3][100] ), .QN(n1137) );
  DFFRX1 \CACHE_reg[3][99]  ( .D(n2376), .CK(clk), .RN(n3781), .Q(
        \CACHE[3][99] ), .QN(n1136) );
  DFFRX1 \CACHE_reg[3][98]  ( .D(n2375), .CK(clk), .RN(n3780), .Q(
        \CACHE[3][98] ), .QN(n1135) );
  DFFRX1 \CACHE_reg[3][97]  ( .D(n2374), .CK(clk), .RN(n3780), .Q(
        \CACHE[3][97] ), .QN(n1134) );
  DFFRX1 \CACHE_reg[3][96]  ( .D(n2373), .CK(clk), .RN(n3780), .Q(
        \CACHE[3][96] ), .QN(n1133) );
  DFFRX1 \CACHE_reg[3][95]  ( .D(n2372), .CK(clk), .RN(n3780), .Q(
        \CACHE[3][95] ), .QN(n1132) );
  DFFRX1 \CACHE_reg[3][94]  ( .D(n2371), .CK(clk), .RN(n3780), .Q(
        \CACHE[3][94] ), .QN(n1131) );
  DFFRX1 \CACHE_reg[3][93]  ( .D(n2370), .CK(clk), .RN(n3780), .Q(
        \CACHE[3][93] ), .QN(n1130) );
  DFFRX1 \CACHE_reg[3][92]  ( .D(n2369), .CK(clk), .RN(n3780), .Q(
        \CACHE[3][92] ), .QN(n1129) );
  DFFRX1 \CACHE_reg[3][91]  ( .D(n2368), .CK(clk), .RN(n3780), .Q(
        \CACHE[3][91] ), .QN(n1128) );
  DFFRX1 \CACHE_reg[3][90]  ( .D(n2367), .CK(clk), .RN(n3780), .Q(
        \CACHE[3][90] ), .QN(n1127) );
  DFFRX1 \CACHE_reg[3][89]  ( .D(n2366), .CK(clk), .RN(n3780), .Q(
        \CACHE[3][89] ), .QN(n1126) );
  DFFRX1 \CACHE_reg[3][88]  ( .D(n2365), .CK(clk), .RN(n3780), .Q(
        \CACHE[3][88] ), .QN(n1125) );
  DFFRX1 \CACHE_reg[3][87]  ( .D(n2364), .CK(clk), .RN(n3780), .Q(
        \CACHE[3][87] ), .QN(n1124) );
  DFFRX1 \CACHE_reg[3][86]  ( .D(n2363), .CK(clk), .RN(n3779), .Q(
        \CACHE[3][86] ), .QN(n1123) );
  DFFRX1 \CACHE_reg[3][85]  ( .D(n2362), .CK(clk), .RN(n3779), .Q(
        \CACHE[3][85] ), .QN(n1122) );
  DFFRX1 \CACHE_reg[3][84]  ( .D(n2361), .CK(clk), .RN(n3779), .Q(
        \CACHE[3][84] ), .QN(n1121) );
  DFFRX1 \CACHE_reg[3][83]  ( .D(n2360), .CK(clk), .RN(n3779), .Q(
        \CACHE[3][83] ), .QN(n1120) );
  DFFRX1 \CACHE_reg[3][82]  ( .D(n2359), .CK(clk), .RN(n3779), .Q(
        \CACHE[3][82] ), .QN(n1119) );
  DFFRX1 \CACHE_reg[3][81]  ( .D(n2358), .CK(clk), .RN(n3779), .Q(
        \CACHE[3][81] ), .QN(n1118) );
  DFFRX1 \CACHE_reg[3][80]  ( .D(n2357), .CK(clk), .RN(n3779), .Q(
        \CACHE[3][80] ), .QN(n1117) );
  DFFRX1 \CACHE_reg[3][79]  ( .D(n2356), .CK(clk), .RN(n3779), .Q(
        \CACHE[3][79] ), .QN(n1116) );
  DFFRX1 \CACHE_reg[3][78]  ( .D(n2355), .CK(clk), .RN(n3779), .Q(
        \CACHE[3][78] ), .QN(n1115) );
  DFFRX1 \CACHE_reg[3][77]  ( .D(n2354), .CK(clk), .RN(n3779), .Q(
        \CACHE[3][77] ), .QN(n1114) );
  DFFRX1 \CACHE_reg[3][76]  ( .D(n2353), .CK(clk), .RN(n3779), .Q(
        \CACHE[3][76] ), .QN(n1113) );
  DFFRX1 \CACHE_reg[3][75]  ( .D(n2352), .CK(clk), .RN(n3779), .Q(
        \CACHE[3][75] ), .QN(n1112) );
  DFFRX1 \CACHE_reg[3][74]  ( .D(n2351), .CK(clk), .RN(n3778), .Q(
        \CACHE[3][74] ), .QN(n1111) );
  DFFRX1 \CACHE_reg[3][73]  ( .D(n2350), .CK(clk), .RN(n3778), .Q(
        \CACHE[3][73] ), .QN(n1110) );
  DFFRX1 \CACHE_reg[3][72]  ( .D(n2349), .CK(clk), .RN(n3778), .Q(
        \CACHE[3][72] ), .QN(n1109) );
  DFFRX1 \CACHE_reg[3][71]  ( .D(n2348), .CK(clk), .RN(n3778), .Q(
        \CACHE[3][71] ), .QN(n1108) );
  DFFRX1 \CACHE_reg[3][70]  ( .D(n2347), .CK(clk), .RN(n3778), .Q(
        \CACHE[3][70] ), .QN(n1107) );
  DFFRX1 \CACHE_reg[3][69]  ( .D(n2346), .CK(clk), .RN(n3778), .Q(
        \CACHE[3][69] ), .QN(n1106) );
  DFFRX1 \CACHE_reg[3][68]  ( .D(n2345), .CK(clk), .RN(n3778), .Q(
        \CACHE[3][68] ), .QN(n1105) );
  DFFRX1 \CACHE_reg[3][67]  ( .D(n2344), .CK(clk), .RN(n3778), .Q(
        \CACHE[3][67] ), .QN(n1104) );
  DFFRX1 \CACHE_reg[3][66]  ( .D(n2343), .CK(clk), .RN(n3778), .Q(
        \CACHE[3][66] ), .QN(n1103) );
  DFFRX1 \CACHE_reg[3][65]  ( .D(n2342), .CK(clk), .RN(n3778), .Q(
        \CACHE[3][65] ), .QN(n1102) );
  DFFRX1 \CACHE_reg[3][64]  ( .D(n2341), .CK(clk), .RN(n3778), .Q(
        \CACHE[3][64] ), .QN(n1101) );
  DFFRX1 \CACHE_reg[3][63]  ( .D(n2340), .CK(clk), .RN(n3778), .Q(
        \CACHE[3][63] ), .QN(n1100) );
  DFFRX1 \CACHE_reg[3][62]  ( .D(n2339), .CK(clk), .RN(n3777), .Q(
        \CACHE[3][62] ), .QN(n1099) );
  DFFRX1 \CACHE_reg[3][61]  ( .D(n2338), .CK(clk), .RN(n3777), .Q(
        \CACHE[3][61] ), .QN(n1098) );
  DFFRX1 \CACHE_reg[3][60]  ( .D(n2337), .CK(clk), .RN(n3777), .Q(
        \CACHE[3][60] ), .QN(n1097) );
  DFFRX1 \CACHE_reg[3][59]  ( .D(n2336), .CK(clk), .RN(n3777), .Q(
        \CACHE[3][59] ), .QN(n1096) );
  DFFRX1 \CACHE_reg[3][58]  ( .D(n2335), .CK(clk), .RN(n3777), .Q(
        \CACHE[3][58] ), .QN(n1095) );
  DFFRX1 \CACHE_reg[3][57]  ( .D(n2334), .CK(clk), .RN(n3777), .Q(
        \CACHE[3][57] ), .QN(n1094) );
  DFFRX1 \CACHE_reg[3][56]  ( .D(n2333), .CK(clk), .RN(n3777), .Q(
        \CACHE[3][56] ), .QN(n1093) );
  DFFRX1 \CACHE_reg[3][55]  ( .D(n2332), .CK(clk), .RN(n3777), .Q(
        \CACHE[3][55] ), .QN(n1092) );
  DFFRX1 \CACHE_reg[3][54]  ( .D(n2331), .CK(clk), .RN(n3777), .Q(
        \CACHE[3][54] ), .QN(n1091) );
  DFFRX1 \CACHE_reg[3][53]  ( .D(n2330), .CK(clk), .RN(n3777), .Q(
        \CACHE[3][53] ), .QN(n1090) );
  DFFRX1 \CACHE_reg[3][52]  ( .D(n2329), .CK(clk), .RN(n3777), .Q(
        \CACHE[3][52] ), .QN(n1089) );
  DFFRX1 \CACHE_reg[3][51]  ( .D(n2328), .CK(clk), .RN(n3777), .Q(
        \CACHE[3][51] ), .QN(n1088) );
  DFFRX1 \CACHE_reg[3][50]  ( .D(n2327), .CK(clk), .RN(n3776), .Q(
        \CACHE[3][50] ), .QN(n1087) );
  DFFRX1 \CACHE_reg[3][49]  ( .D(n2326), .CK(clk), .RN(n3776), .Q(
        \CACHE[3][49] ), .QN(n1086) );
  DFFRX1 \CACHE_reg[3][48]  ( .D(n2325), .CK(clk), .RN(n3776), .Q(
        \CACHE[3][48] ), .QN(n1085) );
  DFFRX1 \CACHE_reg[3][47]  ( .D(n2324), .CK(clk), .RN(n3776), .Q(
        \CACHE[3][47] ), .QN(n1084) );
  DFFRX1 \CACHE_reg[3][46]  ( .D(n2323), .CK(clk), .RN(n3776), .Q(
        \CACHE[3][46] ), .QN(n1083) );
  DFFRX1 \CACHE_reg[3][45]  ( .D(n2322), .CK(clk), .RN(n3776), .Q(
        \CACHE[3][45] ), .QN(n1082) );
  DFFRX1 \CACHE_reg[3][44]  ( .D(n2321), .CK(clk), .RN(n3776), .Q(
        \CACHE[3][44] ), .QN(n1081) );
  DFFRX1 \CACHE_reg[3][43]  ( .D(n2320), .CK(clk), .RN(n3776), .Q(
        \CACHE[3][43] ), .QN(n1080) );
  DFFRX1 \CACHE_reg[3][42]  ( .D(n2319), .CK(clk), .RN(n3776), .Q(
        \CACHE[3][42] ), .QN(n1079) );
  DFFRX1 \CACHE_reg[3][41]  ( .D(n2318), .CK(clk), .RN(n3776), .Q(
        \CACHE[3][41] ), .QN(n1078) );
  DFFRX1 \CACHE_reg[3][40]  ( .D(n2317), .CK(clk), .RN(n3776), .Q(
        \CACHE[3][40] ), .QN(n1077) );
  DFFRX1 \CACHE_reg[3][39]  ( .D(n2316), .CK(clk), .RN(n3776), .Q(
        \CACHE[3][39] ), .QN(n1076) );
  DFFRX1 \CACHE_reg[3][38]  ( .D(n2315), .CK(clk), .RN(n3775), .Q(
        \CACHE[3][38] ), .QN(n1075) );
  DFFRX1 \CACHE_reg[3][37]  ( .D(n2314), .CK(clk), .RN(n3775), .Q(
        \CACHE[3][37] ), .QN(n1074) );
  DFFRX1 \CACHE_reg[3][36]  ( .D(n2313), .CK(clk), .RN(n3775), .Q(
        \CACHE[3][36] ), .QN(n1073) );
  DFFRX1 \CACHE_reg[3][35]  ( .D(n2312), .CK(clk), .RN(n3775), .Q(
        \CACHE[3][35] ), .QN(n1072) );
  DFFRX1 \CACHE_reg[3][34]  ( .D(n2311), .CK(clk), .RN(n3775), .Q(
        \CACHE[3][34] ), .QN(n1071) );
  DFFRX1 \CACHE_reg[3][33]  ( .D(n2310), .CK(clk), .RN(n3775), .Q(
        \CACHE[3][33] ), .QN(n1070) );
  DFFRX1 \CACHE_reg[3][32]  ( .D(n2309), .CK(clk), .RN(n3775), .Q(
        \CACHE[3][32] ), .QN(n1069) );
  DFFRX1 \CACHE_reg[3][31]  ( .D(n2308), .CK(clk), .RN(n3775), .Q(
        \CACHE[3][31] ), .QN(n1068) );
  DFFRX1 \CACHE_reg[3][30]  ( .D(n2307), .CK(clk), .RN(n3775), .Q(
        \CACHE[3][30] ), .QN(n1067) );
  DFFRX1 \CACHE_reg[3][29]  ( .D(n2306), .CK(clk), .RN(n3775), .Q(
        \CACHE[3][29] ), .QN(n1066) );
  DFFRX1 \CACHE_reg[3][28]  ( .D(n2305), .CK(clk), .RN(n3775), .Q(
        \CACHE[3][28] ), .QN(n1065) );
  DFFRX1 \CACHE_reg[3][27]  ( .D(n2304), .CK(clk), .RN(n3775), .Q(
        \CACHE[3][27] ), .QN(n1064) );
  DFFRX1 \CACHE_reg[3][26]  ( .D(n2303), .CK(clk), .RN(n3774), .Q(
        \CACHE[3][26] ), .QN(n1063) );
  DFFRX1 \CACHE_reg[3][25]  ( .D(n2302), .CK(clk), .RN(n3774), .Q(
        \CACHE[3][25] ), .QN(n1062) );
  DFFRX1 \CACHE_reg[3][24]  ( .D(n2301), .CK(clk), .RN(n3774), .Q(
        \CACHE[3][24] ), .QN(n1061) );
  DFFRX1 \CACHE_reg[3][23]  ( .D(n2300), .CK(clk), .RN(n3774), .Q(
        \CACHE[3][23] ), .QN(n1060) );
  DFFRX1 \CACHE_reg[3][22]  ( .D(n2299), .CK(clk), .RN(n3774), .Q(
        \CACHE[3][22] ), .QN(n1059) );
  DFFRX1 \CACHE_reg[3][21]  ( .D(n2298), .CK(clk), .RN(n3774), .Q(
        \CACHE[3][21] ), .QN(n1058) );
  DFFRX1 \CACHE_reg[3][20]  ( .D(n2297), .CK(clk), .RN(n3774), .Q(
        \CACHE[3][20] ), .QN(n1057) );
  DFFRX1 \CACHE_reg[3][19]  ( .D(n2296), .CK(clk), .RN(n3774), .Q(
        \CACHE[3][19] ), .QN(n1056) );
  DFFRX1 \CACHE_reg[3][18]  ( .D(n2295), .CK(clk), .RN(n3774), .Q(
        \CACHE[3][18] ), .QN(n1055) );
  DFFRX1 \CACHE_reg[3][17]  ( .D(n2294), .CK(clk), .RN(n3774), .Q(
        \CACHE[3][17] ), .QN(n1054) );
  DFFRX1 \CACHE_reg[3][16]  ( .D(n2293), .CK(clk), .RN(n3774), .Q(
        \CACHE[3][16] ), .QN(n1053) );
  DFFRX1 \CACHE_reg[3][15]  ( .D(n2292), .CK(clk), .RN(n3774), .Q(
        \CACHE[3][15] ), .QN(n1052) );
  DFFRX1 \CACHE_reg[3][14]  ( .D(n2291), .CK(clk), .RN(n3773), .Q(
        \CACHE[3][14] ), .QN(n1051) );
  DFFRX1 \CACHE_reg[3][13]  ( .D(n2290), .CK(clk), .RN(n3773), .Q(
        \CACHE[3][13] ), .QN(n1050) );
  DFFRX1 \CACHE_reg[3][12]  ( .D(n2289), .CK(clk), .RN(n3773), .Q(
        \CACHE[3][12] ), .QN(n1049) );
  DFFRX1 \CACHE_reg[3][11]  ( .D(n2288), .CK(clk), .RN(n3773), .Q(
        \CACHE[3][11] ), .QN(n1048) );
  DFFRX1 \CACHE_reg[3][10]  ( .D(n2287), .CK(clk), .RN(n3773), .Q(
        \CACHE[3][10] ), .QN(n1047) );
  DFFRX1 \CACHE_reg[3][9]  ( .D(n2286), .CK(clk), .RN(n3773), .Q(\CACHE[3][9] ), .QN(n1046) );
  DFFRX1 \CACHE_reg[3][8]  ( .D(n2285), .CK(clk), .RN(n3773), .Q(\CACHE[3][8] ), .QN(n1045) );
  DFFRX1 \CACHE_reg[3][7]  ( .D(n2284), .CK(clk), .RN(n3773), .Q(\CACHE[3][7] ), .QN(n1044) );
  DFFRX1 \CACHE_reg[3][6]  ( .D(n2283), .CK(clk), .RN(n3773), .Q(\CACHE[3][6] ), .QN(n1043) );
  DFFRX1 \CACHE_reg[3][5]  ( .D(n2282), .CK(clk), .RN(n3773), .Q(\CACHE[3][5] ), .QN(n1042) );
  DFFRX1 \CACHE_reg[3][4]  ( .D(n2281), .CK(clk), .RN(n3773), .Q(\CACHE[3][4] ), .QN(n1041) );
  DFFRX1 \CACHE_reg[3][3]  ( .D(n2280), .CK(clk), .RN(n3773), .Q(\CACHE[3][3] ), .QN(n1040) );
  DFFRX1 \CACHE_reg[3][2]  ( .D(n2279), .CK(clk), .RN(n3772), .Q(\CACHE[3][2] ), .QN(n1039) );
  DFFRX1 \CACHE_reg[3][1]  ( .D(n2278), .CK(clk), .RN(n3772), .Q(\CACHE[3][1] ), .QN(n1038) );
  DFFRX1 \CACHE_reg[3][0]  ( .D(n2277), .CK(clk), .RN(n3772), .Q(\CACHE[3][0] ), .QN(n1037) );
  DFFRX1 \CACHE_reg[5][118]  ( .D(n2705), .CK(clk), .RN(n3808), .Q(
        \CACHE[5][118] ), .QN(n1465) );
  DFFRX1 \CACHE_reg[5][117]  ( .D(n2704), .CK(clk), .RN(n3808), .Q(
        \CACHE[5][117] ), .QN(n1464) );
  DFFRX1 \CACHE_reg[5][116]  ( .D(n2703), .CK(clk), .RN(n3808), .Q(
        \CACHE[5][116] ), .QN(n1463) );
  DFFRX1 \CACHE_reg[5][115]  ( .D(n2702), .CK(clk), .RN(n3808), .Q(
        \CACHE[5][115] ), .QN(n1462) );
  DFFRX1 \CACHE_reg[5][114]  ( .D(n2701), .CK(clk), .RN(n3808), .Q(
        \CACHE[5][114] ), .QN(n1461) );
  DFFRX1 \CACHE_reg[5][113]  ( .D(n2700), .CK(clk), .RN(n3808), .Q(
        \CACHE[5][113] ), .QN(n1460) );
  DFFRX1 \CACHE_reg[5][112]  ( .D(n2699), .CK(clk), .RN(n3807), .Q(
        \CACHE[5][112] ), .QN(n1459) );
  DFFRX1 \CACHE_reg[5][111]  ( .D(n2698), .CK(clk), .RN(n3807), .Q(
        \CACHE[5][111] ), .QN(n1458) );
  DFFRX1 \CACHE_reg[5][110]  ( .D(n2697), .CK(clk), .RN(n3807), .Q(
        \CACHE[5][110] ), .QN(n1457) );
  DFFRX1 \CACHE_reg[5][109]  ( .D(n2696), .CK(clk), .RN(n3807), .Q(
        \CACHE[5][109] ), .QN(n1456) );
  DFFRX1 \CACHE_reg[5][108]  ( .D(n2695), .CK(clk), .RN(n3807), .Q(
        \CACHE[5][108] ), .QN(n1455) );
  DFFRX1 \CACHE_reg[5][107]  ( .D(n2694), .CK(clk), .RN(n3807), .Q(
        \CACHE[5][107] ), .QN(n1454) );
  DFFRX1 \CACHE_reg[5][106]  ( .D(n2693), .CK(clk), .RN(n3807), .Q(
        \CACHE[5][106] ), .QN(n1453) );
  DFFRX1 \CACHE_reg[5][105]  ( .D(n2692), .CK(clk), .RN(n3807), .Q(
        \CACHE[5][105] ), .QN(n1452) );
  DFFRX1 \CACHE_reg[5][104]  ( .D(n2691), .CK(clk), .RN(n3807), .Q(
        \CACHE[5][104] ), .QN(n1451) );
  DFFRX1 \CACHE_reg[5][103]  ( .D(n2690), .CK(clk), .RN(n3807), .Q(
        \CACHE[5][103] ), .QN(n1450) );
  DFFRX1 \CACHE_reg[5][102]  ( .D(n2689), .CK(clk), .RN(n3807), .Q(
        \CACHE[5][102] ), .QN(n1449) );
  DFFRX1 \CACHE_reg[5][101]  ( .D(n2688), .CK(clk), .RN(n3807), .Q(
        \CACHE[5][101] ), .QN(n1448) );
  DFFRX1 \CACHE_reg[5][100]  ( .D(n2687), .CK(clk), .RN(n3806), .Q(
        \CACHE[5][100] ), .QN(n1447) );
  DFFRX1 \CACHE_reg[5][99]  ( .D(n2686), .CK(clk), .RN(n3806), .Q(
        \CACHE[5][99] ), .QN(n1446) );
  DFFRX1 \CACHE_reg[5][98]  ( .D(n2685), .CK(clk), .RN(n3806), .Q(
        \CACHE[5][98] ), .QN(n1445) );
  DFFRX1 \CACHE_reg[5][97]  ( .D(n2684), .CK(clk), .RN(n3806), .Q(
        \CACHE[5][97] ), .QN(n1444) );
  DFFRX1 \CACHE_reg[5][96]  ( .D(n2683), .CK(clk), .RN(n3806), .Q(
        \CACHE[5][96] ), .QN(n1443) );
  DFFRX1 \CACHE_reg[5][95]  ( .D(n2682), .CK(clk), .RN(n3806), .Q(
        \CACHE[5][95] ), .QN(n1442) );
  DFFRX1 \CACHE_reg[5][94]  ( .D(n2681), .CK(clk), .RN(n3806), .Q(
        \CACHE[5][94] ), .QN(n1441) );
  DFFRX1 \CACHE_reg[5][93]  ( .D(n2680), .CK(clk), .RN(n3806), .Q(
        \CACHE[5][93] ), .QN(n1440) );
  DFFRX1 \CACHE_reg[5][92]  ( .D(n2679), .CK(clk), .RN(n3806), .Q(
        \CACHE[5][92] ), .QN(n1439) );
  DFFRX1 \CACHE_reg[5][91]  ( .D(n2678), .CK(clk), .RN(n3806), .Q(
        \CACHE[5][91] ), .QN(n1438) );
  DFFRX1 \CACHE_reg[5][90]  ( .D(n2677), .CK(clk), .RN(n3806), .Q(
        \CACHE[5][90] ), .QN(n1437) );
  DFFRX1 \CACHE_reg[5][89]  ( .D(n2676), .CK(clk), .RN(n3806), .Q(
        \CACHE[5][89] ), .QN(n1436) );
  DFFRX1 \CACHE_reg[5][88]  ( .D(n2675), .CK(clk), .RN(n3805), .Q(
        \CACHE[5][88] ), .QN(n1435) );
  DFFRX1 \CACHE_reg[5][87]  ( .D(n2674), .CK(clk), .RN(n3805), .Q(
        \CACHE[5][87] ), .QN(n1434) );
  DFFRX1 \CACHE_reg[5][86]  ( .D(n2673), .CK(clk), .RN(n3805), .Q(
        \CACHE[5][86] ), .QN(n1433) );
  DFFRX1 \CACHE_reg[5][85]  ( .D(n2672), .CK(clk), .RN(n3805), .Q(
        \CACHE[5][85] ), .QN(n1432) );
  DFFRX1 \CACHE_reg[5][84]  ( .D(n2671), .CK(clk), .RN(n3805), .Q(
        \CACHE[5][84] ), .QN(n1431) );
  DFFRX1 \CACHE_reg[5][83]  ( .D(n2670), .CK(clk), .RN(n3805), .Q(
        \CACHE[5][83] ), .QN(n1430) );
  DFFRX1 \CACHE_reg[5][82]  ( .D(n2669), .CK(clk), .RN(n3805), .Q(
        \CACHE[5][82] ), .QN(n1429) );
  DFFRX1 \CACHE_reg[5][81]  ( .D(n2668), .CK(clk), .RN(n3805), .Q(
        \CACHE[5][81] ), .QN(n1428) );
  DFFRX1 \CACHE_reg[5][80]  ( .D(n2667), .CK(clk), .RN(n3805), .Q(
        \CACHE[5][80] ), .QN(n1427) );
  DFFRX1 \CACHE_reg[5][79]  ( .D(n2666), .CK(clk), .RN(n3805), .Q(
        \CACHE[5][79] ), .QN(n1426) );
  DFFRX1 \CACHE_reg[5][78]  ( .D(n2665), .CK(clk), .RN(n3805), .Q(
        \CACHE[5][78] ), .QN(n1425) );
  DFFRX1 \CACHE_reg[5][77]  ( .D(n2664), .CK(clk), .RN(n3805), .Q(
        \CACHE[5][77] ), .QN(n1424) );
  DFFRX1 \CACHE_reg[5][76]  ( .D(n2663), .CK(clk), .RN(n3804), .Q(
        \CACHE[5][76] ), .QN(n1423) );
  DFFRX1 \CACHE_reg[5][75]  ( .D(n2662), .CK(clk), .RN(n3804), .Q(
        \CACHE[5][75] ), .QN(n1422) );
  DFFRX1 \CACHE_reg[5][74]  ( .D(n2661), .CK(clk), .RN(n3804), .Q(
        \CACHE[5][74] ), .QN(n1421) );
  DFFRX1 \CACHE_reg[5][73]  ( .D(n2660), .CK(clk), .RN(n3804), .Q(
        \CACHE[5][73] ), .QN(n1420) );
  DFFRX1 \CACHE_reg[5][72]  ( .D(n2659), .CK(clk), .RN(n3804), .Q(
        \CACHE[5][72] ), .QN(n1419) );
  DFFRX1 \CACHE_reg[5][71]  ( .D(n2658), .CK(clk), .RN(n3804), .Q(
        \CACHE[5][71] ), .QN(n1418) );
  DFFRX1 \CACHE_reg[5][70]  ( .D(n2657), .CK(clk), .RN(n3804), .Q(
        \CACHE[5][70] ), .QN(n1417) );
  DFFRX1 \CACHE_reg[5][69]  ( .D(n2656), .CK(clk), .RN(n3804), .Q(
        \CACHE[5][69] ), .QN(n1416) );
  DFFRX1 \CACHE_reg[5][68]  ( .D(n2655), .CK(clk), .RN(n3804), .Q(
        \CACHE[5][68] ), .QN(n1415) );
  DFFRX1 \CACHE_reg[5][67]  ( .D(n2654), .CK(clk), .RN(n3804), .Q(
        \CACHE[5][67] ), .QN(n1414) );
  DFFRX1 \CACHE_reg[5][66]  ( .D(n2653), .CK(clk), .RN(n3804), .Q(
        \CACHE[5][66] ), .QN(n1413) );
  DFFRX1 \CACHE_reg[5][65]  ( .D(n2652), .CK(clk), .RN(n3804), .Q(
        \CACHE[5][65] ), .QN(n1412) );
  DFFRX1 \CACHE_reg[5][64]  ( .D(n2651), .CK(clk), .RN(n3803), .Q(
        \CACHE[5][64] ), .QN(n1411) );
  DFFRX1 \CACHE_reg[5][63]  ( .D(n2650), .CK(clk), .RN(n3803), .Q(
        \CACHE[5][63] ), .QN(n1410) );
  DFFRX1 \CACHE_reg[5][62]  ( .D(n2649), .CK(clk), .RN(n3803), .Q(
        \CACHE[5][62] ), .QN(n1409) );
  DFFRX1 \CACHE_reg[5][61]  ( .D(n2648), .CK(clk), .RN(n3803), .Q(
        \CACHE[5][61] ), .QN(n1408) );
  DFFRX1 \CACHE_reg[5][60]  ( .D(n2647), .CK(clk), .RN(n3803), .Q(
        \CACHE[5][60] ), .QN(n1407) );
  DFFRX1 \CACHE_reg[5][59]  ( .D(n2646), .CK(clk), .RN(n3803), .Q(
        \CACHE[5][59] ), .QN(n1406) );
  DFFRX1 \CACHE_reg[5][58]  ( .D(n2645), .CK(clk), .RN(n3803), .Q(
        \CACHE[5][58] ), .QN(n1405) );
  DFFRX1 \CACHE_reg[5][57]  ( .D(n2644), .CK(clk), .RN(n3803), .Q(
        \CACHE[5][57] ), .QN(n1404) );
  DFFRX1 \CACHE_reg[5][56]  ( .D(n2643), .CK(clk), .RN(n3803), .Q(
        \CACHE[5][56] ), .QN(n1403) );
  DFFRX1 \CACHE_reg[5][55]  ( .D(n2642), .CK(clk), .RN(n3803), .Q(
        \CACHE[5][55] ), .QN(n1402) );
  DFFRX1 \CACHE_reg[5][54]  ( .D(n2641), .CK(clk), .RN(n3803), .Q(
        \CACHE[5][54] ), .QN(n1401) );
  DFFRX1 \CACHE_reg[5][53]  ( .D(n2640), .CK(clk), .RN(n3803), .Q(
        \CACHE[5][53] ), .QN(n1400) );
  DFFRX1 \CACHE_reg[5][52]  ( .D(n2639), .CK(clk), .RN(n3802), .Q(
        \CACHE[5][52] ), .QN(n1399) );
  DFFRX1 \CACHE_reg[5][51]  ( .D(n2638), .CK(clk), .RN(n3802), .Q(
        \CACHE[5][51] ), .QN(n1398) );
  DFFRX1 \CACHE_reg[5][50]  ( .D(n2637), .CK(clk), .RN(n3802), .Q(
        \CACHE[5][50] ), .QN(n1397) );
  DFFRX1 \CACHE_reg[5][49]  ( .D(n2636), .CK(clk), .RN(n3802), .Q(
        \CACHE[5][49] ), .QN(n1396) );
  DFFRX1 \CACHE_reg[5][48]  ( .D(n2635), .CK(clk), .RN(n3802), .Q(
        \CACHE[5][48] ), .QN(n1395) );
  DFFRX1 \CACHE_reg[5][47]  ( .D(n2634), .CK(clk), .RN(n3802), .Q(
        \CACHE[5][47] ), .QN(n1394) );
  DFFRX1 \CACHE_reg[5][46]  ( .D(n2633), .CK(clk), .RN(n3802), .Q(
        \CACHE[5][46] ), .QN(n1393) );
  DFFRX1 \CACHE_reg[5][45]  ( .D(n2632), .CK(clk), .RN(n3802), .Q(
        \CACHE[5][45] ), .QN(n1392) );
  DFFRX1 \CACHE_reg[5][44]  ( .D(n2631), .CK(clk), .RN(n3802), .Q(
        \CACHE[5][44] ), .QN(n1391) );
  DFFRX1 \CACHE_reg[5][43]  ( .D(n2630), .CK(clk), .RN(n3802), .Q(
        \CACHE[5][43] ), .QN(n1390) );
  DFFRX1 \CACHE_reg[5][42]  ( .D(n2629), .CK(clk), .RN(n3802), .Q(
        \CACHE[5][42] ), .QN(n1389) );
  DFFRX1 \CACHE_reg[5][41]  ( .D(n2628), .CK(clk), .RN(n3802), .Q(
        \CACHE[5][41] ), .QN(n1388) );
  DFFRX1 \CACHE_reg[5][40]  ( .D(n2627), .CK(clk), .RN(n3801), .Q(
        \CACHE[5][40] ), .QN(n1387) );
  DFFRX1 \CACHE_reg[5][39]  ( .D(n2626), .CK(clk), .RN(n3801), .Q(
        \CACHE[5][39] ), .QN(n1386) );
  DFFRX1 \CACHE_reg[5][38]  ( .D(n2625), .CK(clk), .RN(n3801), .Q(
        \CACHE[5][38] ), .QN(n1385) );
  DFFRX1 \CACHE_reg[5][37]  ( .D(n2624), .CK(clk), .RN(n3801), .Q(
        \CACHE[5][37] ), .QN(n1384) );
  DFFRX1 \CACHE_reg[5][36]  ( .D(n2623), .CK(clk), .RN(n3801), .Q(
        \CACHE[5][36] ), .QN(n1383) );
  DFFRX1 \CACHE_reg[5][35]  ( .D(n2622), .CK(clk), .RN(n3801), .Q(
        \CACHE[5][35] ), .QN(n1382) );
  DFFRX1 \CACHE_reg[5][34]  ( .D(n2621), .CK(clk), .RN(n3801), .Q(
        \CACHE[5][34] ), .QN(n1381) );
  DFFRX1 \CACHE_reg[5][33]  ( .D(n2620), .CK(clk), .RN(n3801), .Q(
        \CACHE[5][33] ), .QN(n1380) );
  DFFRX1 \CACHE_reg[5][32]  ( .D(n2619), .CK(clk), .RN(n3801), .Q(
        \CACHE[5][32] ), .QN(n1379) );
  DFFRX1 \CACHE_reg[5][31]  ( .D(n2618), .CK(clk), .RN(n3801), .Q(
        \CACHE[5][31] ), .QN(n1378) );
  DFFRX1 \CACHE_reg[5][30]  ( .D(n2617), .CK(clk), .RN(n3801), .Q(
        \CACHE[5][30] ), .QN(n1377) );
  DFFRX1 \CACHE_reg[5][29]  ( .D(n2616), .CK(clk), .RN(n3801), .Q(
        \CACHE[5][29] ), .QN(n1376) );
  DFFRX1 \CACHE_reg[5][28]  ( .D(n2615), .CK(clk), .RN(n3800), .Q(
        \CACHE[5][28] ), .QN(n1375) );
  DFFRX1 \CACHE_reg[5][27]  ( .D(n2614), .CK(clk), .RN(n3800), .Q(
        \CACHE[5][27] ), .QN(n1374) );
  DFFRX1 \CACHE_reg[5][26]  ( .D(n2613), .CK(clk), .RN(n3800), .Q(
        \CACHE[5][26] ), .QN(n1373) );
  DFFRX1 \CACHE_reg[5][25]  ( .D(n2612), .CK(clk), .RN(n3800), .Q(
        \CACHE[5][25] ), .QN(n1372) );
  DFFRX1 \CACHE_reg[5][24]  ( .D(n2611), .CK(clk), .RN(n3800), .Q(
        \CACHE[5][24] ), .QN(n1371) );
  DFFRX1 \CACHE_reg[5][23]  ( .D(n2610), .CK(clk), .RN(n3800), .Q(
        \CACHE[5][23] ), .QN(n1370) );
  DFFRX1 \CACHE_reg[5][22]  ( .D(n2609), .CK(clk), .RN(n3800), .Q(
        \CACHE[5][22] ), .QN(n1369) );
  DFFRX1 \CACHE_reg[5][21]  ( .D(n2608), .CK(clk), .RN(n3800), .Q(
        \CACHE[5][21] ), .QN(n1368) );
  DFFRX1 \CACHE_reg[5][20]  ( .D(n2607), .CK(clk), .RN(n3800), .Q(
        \CACHE[5][20] ), .QN(n1367) );
  DFFRX1 \CACHE_reg[5][19]  ( .D(n2606), .CK(clk), .RN(n3800), .Q(
        \CACHE[5][19] ), .QN(n1366) );
  DFFRX1 \CACHE_reg[5][18]  ( .D(n2605), .CK(clk), .RN(n3800), .Q(
        \CACHE[5][18] ), .QN(n1365) );
  DFFRX1 \CACHE_reg[5][17]  ( .D(n2604), .CK(clk), .RN(n3800), .Q(
        \CACHE[5][17] ), .QN(n1364) );
  DFFRX1 \CACHE_reg[5][16]  ( .D(n2603), .CK(clk), .RN(n3799), .Q(
        \CACHE[5][16] ), .QN(n1363) );
  DFFRX1 \CACHE_reg[5][15]  ( .D(n2602), .CK(clk), .RN(n3799), .Q(
        \CACHE[5][15] ), .QN(n1362) );
  DFFRX1 \CACHE_reg[5][14]  ( .D(n2601), .CK(clk), .RN(n3799), .Q(
        \CACHE[5][14] ), .QN(n1361) );
  DFFRX1 \CACHE_reg[5][13]  ( .D(n2600), .CK(clk), .RN(n3799), .Q(
        \CACHE[5][13] ), .QN(n1360) );
  DFFRX1 \CACHE_reg[5][12]  ( .D(n2599), .CK(clk), .RN(n3799), .Q(
        \CACHE[5][12] ), .QN(n1359) );
  DFFRX1 \CACHE_reg[5][11]  ( .D(n2598), .CK(clk), .RN(n3799), .Q(
        \CACHE[5][11] ), .QN(n1358) );
  DFFRX1 \CACHE_reg[5][10]  ( .D(n2597), .CK(clk), .RN(n3799), .Q(
        \CACHE[5][10] ), .QN(n1357) );
  DFFRX1 \CACHE_reg[5][9]  ( .D(n2596), .CK(clk), .RN(n3799), .Q(\CACHE[5][9] ), .QN(n1356) );
  DFFRX1 \CACHE_reg[5][8]  ( .D(n2595), .CK(clk), .RN(n3799), .Q(\CACHE[5][8] ), .QN(n1355) );
  DFFRX1 \CACHE_reg[5][7]  ( .D(n2594), .CK(clk), .RN(n3799), .Q(\CACHE[5][7] ), .QN(n1354) );
  DFFRX1 \CACHE_reg[5][6]  ( .D(n2593), .CK(clk), .RN(n3799), .Q(\CACHE[5][6] ), .QN(n1353) );
  DFFRX1 \CACHE_reg[5][5]  ( .D(n2592), .CK(clk), .RN(n3799), .Q(\CACHE[5][5] ), .QN(n1352) );
  DFFRX1 \CACHE_reg[5][4]  ( .D(n2591), .CK(clk), .RN(n3798), .Q(\CACHE[5][4] ), .QN(n1351) );
  DFFRX1 \CACHE_reg[5][3]  ( .D(n2590), .CK(clk), .RN(n3798), .Q(\CACHE[5][3] ), .QN(n1350) );
  DFFRX1 \CACHE_reg[5][2]  ( .D(n2589), .CK(clk), .RN(n3798), .Q(\CACHE[5][2] ), .QN(n1349) );
  DFFRX1 \CACHE_reg[5][1]  ( .D(n2588), .CK(clk), .RN(n3798), .Q(\CACHE[5][1] ), .QN(n1348) );
  DFFRX1 \CACHE_reg[5][0]  ( .D(n2587), .CK(clk), .RN(n3798), .Q(\CACHE[5][0] ), .QN(n1347) );
  DFFRX1 \CACHE_reg[1][118]  ( .D(n2085), .CK(clk), .RN(n3756), .Q(
        \CACHE[1][118] ), .QN(n845) );
  DFFRX1 \CACHE_reg[1][117]  ( .D(n2084), .CK(clk), .RN(n3756), .Q(
        \CACHE[1][117] ), .QN(n844) );
  DFFRX1 \CACHE_reg[1][116]  ( .D(n2083), .CK(clk), .RN(n3756), .Q(
        \CACHE[1][116] ), .QN(n843) );
  DFFRX1 \CACHE_reg[1][115]  ( .D(n2082), .CK(clk), .RN(n3756), .Q(
        \CACHE[1][115] ), .QN(n842) );
  DFFRX1 \CACHE_reg[1][114]  ( .D(n2081), .CK(clk), .RN(n3756), .Q(
        \CACHE[1][114] ), .QN(n841) );
  DFFRX1 \CACHE_reg[1][113]  ( .D(n2080), .CK(clk), .RN(n3756), .Q(
        \CACHE[1][113] ), .QN(n840) );
  DFFRX1 \CACHE_reg[1][112]  ( .D(n2079), .CK(clk), .RN(n3756), .Q(
        \CACHE[1][112] ), .QN(n839) );
  DFFRX1 \CACHE_reg[1][111]  ( .D(n2078), .CK(clk), .RN(n3756), .Q(
        \CACHE[1][111] ), .QN(n838) );
  DFFRX1 \CACHE_reg[1][110]  ( .D(n2077), .CK(clk), .RN(n3756), .Q(
        \CACHE[1][110] ), .QN(n837) );
  DFFRX1 \CACHE_reg[1][109]  ( .D(n2076), .CK(clk), .RN(n3756), .Q(
        \CACHE[1][109] ), .QN(n836) );
  DFFRX1 \CACHE_reg[1][108]  ( .D(n2075), .CK(clk), .RN(n3755), .Q(
        \CACHE[1][108] ), .QN(n835) );
  DFFRX1 \CACHE_reg[1][107]  ( .D(n2074), .CK(clk), .RN(n3755), .Q(
        \CACHE[1][107] ), .QN(n834) );
  DFFRX1 \CACHE_reg[1][106]  ( .D(n2073), .CK(clk), .RN(n3755), .Q(
        \CACHE[1][106] ), .QN(n833) );
  DFFRX1 \CACHE_reg[1][105]  ( .D(n2072), .CK(clk), .RN(n3755), .Q(
        \CACHE[1][105] ), .QN(n832) );
  DFFRX1 \CACHE_reg[1][104]  ( .D(n2071), .CK(clk), .RN(n3755), .Q(
        \CACHE[1][104] ), .QN(n831) );
  DFFRX1 \CACHE_reg[1][103]  ( .D(n2070), .CK(clk), .RN(n3755), .Q(
        \CACHE[1][103] ), .QN(n830) );
  DFFRX1 \CACHE_reg[1][102]  ( .D(n2069), .CK(clk), .RN(n3755), .Q(
        \CACHE[1][102] ), .QN(n829) );
  DFFRX1 \CACHE_reg[1][101]  ( .D(n2068), .CK(clk), .RN(n3755), .Q(
        \CACHE[1][101] ), .QN(n828) );
  DFFRX1 \CACHE_reg[1][100]  ( .D(n2067), .CK(clk), .RN(n3755), .Q(
        \CACHE[1][100] ), .QN(n827) );
  DFFRX1 \CACHE_reg[1][99]  ( .D(n2066), .CK(clk), .RN(n3755), .Q(
        \CACHE[1][99] ), .QN(n826) );
  DFFRX1 \CACHE_reg[1][98]  ( .D(n2065), .CK(clk), .RN(n3755), .Q(
        \CACHE[1][98] ), .QN(n825) );
  DFFRX1 \CACHE_reg[1][97]  ( .D(n2064), .CK(clk), .RN(n3755), .Q(
        \CACHE[1][97] ), .QN(n824) );
  DFFRX1 \CACHE_reg[1][96]  ( .D(n2063), .CK(clk), .RN(n3754), .Q(
        \CACHE[1][96] ), .QN(n823) );
  DFFRX1 \CACHE_reg[1][95]  ( .D(n2062), .CK(clk), .RN(n3754), .Q(
        \CACHE[1][95] ), .QN(n822) );
  DFFRX1 \CACHE_reg[1][94]  ( .D(n2061), .CK(clk), .RN(n3754), .Q(
        \CACHE[1][94] ), .QN(n821) );
  DFFRX1 \CACHE_reg[1][93]  ( .D(n2060), .CK(clk), .RN(n3754), .Q(
        \CACHE[1][93] ), .QN(n820) );
  DFFRX1 \CACHE_reg[1][92]  ( .D(n2059), .CK(clk), .RN(n3754), .Q(
        \CACHE[1][92] ), .QN(n819) );
  DFFRX1 \CACHE_reg[1][91]  ( .D(n2058), .CK(clk), .RN(n3754), .Q(
        \CACHE[1][91] ), .QN(n818) );
  DFFRX1 \CACHE_reg[1][90]  ( .D(n2057), .CK(clk), .RN(n3754), .Q(
        \CACHE[1][90] ), .QN(n817) );
  DFFRX1 \CACHE_reg[1][89]  ( .D(n2056), .CK(clk), .RN(n3754), .Q(
        \CACHE[1][89] ), .QN(n816) );
  DFFRX1 \CACHE_reg[1][88]  ( .D(n2055), .CK(clk), .RN(n3754), .Q(
        \CACHE[1][88] ), .QN(n815) );
  DFFRX1 \CACHE_reg[1][87]  ( .D(n2054), .CK(clk), .RN(n3754), .Q(
        \CACHE[1][87] ), .QN(n814) );
  DFFRX1 \CACHE_reg[1][86]  ( .D(n2053), .CK(clk), .RN(n3754), .Q(
        \CACHE[1][86] ), .QN(n813) );
  DFFRX1 \CACHE_reg[1][85]  ( .D(n2052), .CK(clk), .RN(n3754), .Q(
        \CACHE[1][85] ), .QN(n812) );
  DFFRX1 \CACHE_reg[1][84]  ( .D(n2051), .CK(clk), .RN(n3753), .Q(
        \CACHE[1][84] ), .QN(n811) );
  DFFRX1 \CACHE_reg[1][83]  ( .D(n2050), .CK(clk), .RN(n3753), .Q(
        \CACHE[1][83] ), .QN(n810) );
  DFFRX1 \CACHE_reg[1][82]  ( .D(n2049), .CK(clk), .RN(n3753), .Q(
        \CACHE[1][82] ), .QN(n809) );
  DFFRX1 \CACHE_reg[1][81]  ( .D(n2048), .CK(clk), .RN(n3753), .Q(
        \CACHE[1][81] ), .QN(n808) );
  DFFRX1 \CACHE_reg[1][80]  ( .D(n2047), .CK(clk), .RN(n3753), .Q(
        \CACHE[1][80] ), .QN(n807) );
  DFFRX1 \CACHE_reg[1][79]  ( .D(n2046), .CK(clk), .RN(n3753), .Q(
        \CACHE[1][79] ), .QN(n806) );
  DFFRX1 \CACHE_reg[1][78]  ( .D(n2045), .CK(clk), .RN(n3753), .Q(
        \CACHE[1][78] ), .QN(n805) );
  DFFRX1 \CACHE_reg[1][77]  ( .D(n2044), .CK(clk), .RN(n3753), .Q(
        \CACHE[1][77] ), .QN(n804) );
  DFFRX1 \CACHE_reg[1][76]  ( .D(n2043), .CK(clk), .RN(n3753), .Q(
        \CACHE[1][76] ), .QN(n803) );
  DFFRX1 \CACHE_reg[1][75]  ( .D(n2042), .CK(clk), .RN(n3753), .Q(
        \CACHE[1][75] ), .QN(n802) );
  DFFRX1 \CACHE_reg[1][74]  ( .D(n2041), .CK(clk), .RN(n3753), .Q(
        \CACHE[1][74] ), .QN(n801) );
  DFFRX1 \CACHE_reg[1][73]  ( .D(n2040), .CK(clk), .RN(n3753), .Q(
        \CACHE[1][73] ), .QN(n800) );
  DFFRX1 \CACHE_reg[1][72]  ( .D(n2039), .CK(clk), .RN(n3752), .Q(
        \CACHE[1][72] ), .QN(n799) );
  DFFRX1 \CACHE_reg[1][71]  ( .D(n2038), .CK(clk), .RN(n3752), .Q(
        \CACHE[1][71] ), .QN(n798) );
  DFFRX1 \CACHE_reg[1][70]  ( .D(n2037), .CK(clk), .RN(n3752), .Q(
        \CACHE[1][70] ), .QN(n797) );
  DFFRX1 \CACHE_reg[1][69]  ( .D(n2036), .CK(clk), .RN(n3752), .Q(
        \CACHE[1][69] ), .QN(n796) );
  DFFRX1 \CACHE_reg[1][68]  ( .D(n2035), .CK(clk), .RN(n3752), .Q(
        \CACHE[1][68] ), .QN(n795) );
  DFFRX1 \CACHE_reg[1][67]  ( .D(n2034), .CK(clk), .RN(n3752), .Q(
        \CACHE[1][67] ), .QN(n794) );
  DFFRX1 \CACHE_reg[1][66]  ( .D(n2033), .CK(clk), .RN(n3752), .Q(
        \CACHE[1][66] ), .QN(n793) );
  DFFRX1 \CACHE_reg[1][65]  ( .D(n2032), .CK(clk), .RN(n3752), .Q(
        \CACHE[1][65] ), .QN(n792) );
  DFFRX1 \CACHE_reg[1][64]  ( .D(n2031), .CK(clk), .RN(n3752), .Q(
        \CACHE[1][64] ), .QN(n791) );
  DFFRX1 \CACHE_reg[1][63]  ( .D(n2030), .CK(clk), .RN(n3752), .Q(
        \CACHE[1][63] ), .QN(n790) );
  DFFRX1 \CACHE_reg[1][62]  ( .D(n2029), .CK(clk), .RN(n3752), .Q(
        \CACHE[1][62] ), .QN(n789) );
  DFFRX1 \CACHE_reg[1][61]  ( .D(n2028), .CK(clk), .RN(n3752), .Q(
        \CACHE[1][61] ), .QN(n788) );
  DFFRX1 \CACHE_reg[1][60]  ( .D(n2027), .CK(clk), .RN(n3751), .Q(
        \CACHE[1][60] ), .QN(n787) );
  DFFRX1 \CACHE_reg[1][59]  ( .D(n2026), .CK(clk), .RN(n3751), .Q(
        \CACHE[1][59] ), .QN(n786) );
  DFFRX1 \CACHE_reg[1][58]  ( .D(n2025), .CK(clk), .RN(n3751), .Q(
        \CACHE[1][58] ), .QN(n785) );
  DFFRX1 \CACHE_reg[1][57]  ( .D(n2024), .CK(clk), .RN(n3751), .Q(
        \CACHE[1][57] ), .QN(n784) );
  DFFRX1 \CACHE_reg[1][56]  ( .D(n2023), .CK(clk), .RN(n3751), .Q(
        \CACHE[1][56] ), .QN(n783) );
  DFFRX1 \CACHE_reg[1][55]  ( .D(n2022), .CK(clk), .RN(n3751), .Q(
        \CACHE[1][55] ), .QN(n782) );
  DFFRX1 \CACHE_reg[1][54]  ( .D(n2021), .CK(clk), .RN(n3751), .Q(
        \CACHE[1][54] ), .QN(n781) );
  DFFRX1 \CACHE_reg[1][53]  ( .D(n2020), .CK(clk), .RN(n3751), .Q(
        \CACHE[1][53] ), .QN(n780) );
  DFFRX1 \CACHE_reg[1][52]  ( .D(n2019), .CK(clk), .RN(n3751), .Q(
        \CACHE[1][52] ), .QN(n779) );
  DFFRX1 \CACHE_reg[1][51]  ( .D(n2018), .CK(clk), .RN(n3751), .Q(
        \CACHE[1][51] ), .QN(n778) );
  DFFRX1 \CACHE_reg[1][50]  ( .D(n2017), .CK(clk), .RN(n3751), .Q(
        \CACHE[1][50] ), .QN(n777) );
  DFFRX1 \CACHE_reg[1][49]  ( .D(n2016), .CK(clk), .RN(n3751), .Q(
        \CACHE[1][49] ), .QN(n776) );
  DFFRX1 \CACHE_reg[1][48]  ( .D(n2015), .CK(clk), .RN(n3750), .Q(
        \CACHE[1][48] ), .QN(n775) );
  DFFRX1 \CACHE_reg[1][47]  ( .D(n2014), .CK(clk), .RN(n3750), .Q(
        \CACHE[1][47] ), .QN(n774) );
  DFFRX1 \CACHE_reg[1][46]  ( .D(n2013), .CK(clk), .RN(n3750), .Q(
        \CACHE[1][46] ), .QN(n773) );
  DFFRX1 \CACHE_reg[1][45]  ( .D(n2012), .CK(clk), .RN(n3750), .Q(
        \CACHE[1][45] ), .QN(n772) );
  DFFRX1 \CACHE_reg[1][44]  ( .D(n2011), .CK(clk), .RN(n3750), .Q(
        \CACHE[1][44] ), .QN(n771) );
  DFFRX1 \CACHE_reg[1][43]  ( .D(n2010), .CK(clk), .RN(n3750), .Q(
        \CACHE[1][43] ), .QN(n770) );
  DFFRX1 \CACHE_reg[1][42]  ( .D(n2009), .CK(clk), .RN(n3750), .Q(
        \CACHE[1][42] ), .QN(n769) );
  DFFRX1 \CACHE_reg[1][41]  ( .D(n2008), .CK(clk), .RN(n3750), .Q(
        \CACHE[1][41] ), .QN(n768) );
  DFFRX1 \CACHE_reg[1][40]  ( .D(n2007), .CK(clk), .RN(n3750), .Q(
        \CACHE[1][40] ), .QN(n767) );
  DFFRX1 \CACHE_reg[1][39]  ( .D(n2006), .CK(clk), .RN(n3750), .Q(
        \CACHE[1][39] ), .QN(n766) );
  DFFRX1 \CACHE_reg[1][38]  ( .D(n2005), .CK(clk), .RN(n3750), .Q(
        \CACHE[1][38] ), .QN(n765) );
  DFFRX1 \CACHE_reg[1][37]  ( .D(n2004), .CK(clk), .RN(n3750), .Q(
        \CACHE[1][37] ), .QN(n764) );
  DFFRX1 \CACHE_reg[1][36]  ( .D(n2003), .CK(clk), .RN(n3749), .Q(
        \CACHE[1][36] ), .QN(n763) );
  DFFRX1 \CACHE_reg[1][35]  ( .D(n2002), .CK(clk), .RN(n3749), .Q(
        \CACHE[1][35] ), .QN(n762) );
  DFFRX1 \CACHE_reg[1][34]  ( .D(n2001), .CK(clk), .RN(n3749), .Q(
        \CACHE[1][34] ), .QN(n761) );
  DFFRX1 \CACHE_reg[1][33]  ( .D(n2000), .CK(clk), .RN(n3749), .Q(
        \CACHE[1][33] ), .QN(n760) );
  DFFRX1 \CACHE_reg[1][32]  ( .D(n1999), .CK(clk), .RN(n3749), .Q(
        \CACHE[1][32] ), .QN(n759) );
  DFFRX1 \CACHE_reg[1][31]  ( .D(n1998), .CK(clk), .RN(n3749), .Q(
        \CACHE[1][31] ), .QN(n758) );
  DFFRX1 \CACHE_reg[1][30]  ( .D(n1997), .CK(clk), .RN(n3749), .Q(
        \CACHE[1][30] ), .QN(n757) );
  DFFRX1 \CACHE_reg[1][29]  ( .D(n1996), .CK(clk), .RN(n3749), .Q(
        \CACHE[1][29] ), .QN(n756) );
  DFFRX1 \CACHE_reg[1][28]  ( .D(n1995), .CK(clk), .RN(n3749), .Q(
        \CACHE[1][28] ), .QN(n755) );
  DFFRX1 \CACHE_reg[1][27]  ( .D(n1994), .CK(clk), .RN(n3749), .Q(
        \CACHE[1][27] ), .QN(n754) );
  DFFRX1 \CACHE_reg[1][26]  ( .D(n1993), .CK(clk), .RN(n3749), .Q(
        \CACHE[1][26] ), .QN(n753) );
  DFFRX1 \CACHE_reg[1][25]  ( .D(n1992), .CK(clk), .RN(n3749), .Q(
        \CACHE[1][25] ), .QN(n752) );
  DFFRX1 \CACHE_reg[1][24]  ( .D(n1991), .CK(clk), .RN(n3748), .Q(
        \CACHE[1][24] ), .QN(n751) );
  DFFRX1 \CACHE_reg[1][23]  ( .D(n1990), .CK(clk), .RN(n3748), .Q(
        \CACHE[1][23] ), .QN(n750) );
  DFFRX1 \CACHE_reg[1][22]  ( .D(n1989), .CK(clk), .RN(n3748), .Q(
        \CACHE[1][22] ), .QN(n749) );
  DFFRX1 \CACHE_reg[1][21]  ( .D(n1988), .CK(clk), .RN(n3748), .Q(
        \CACHE[1][21] ), .QN(n748) );
  DFFRX1 \CACHE_reg[1][20]  ( .D(n1987), .CK(clk), .RN(n3748), .Q(
        \CACHE[1][20] ), .QN(n747) );
  DFFRX1 \CACHE_reg[1][19]  ( .D(n1986), .CK(clk), .RN(n3748), .Q(
        \CACHE[1][19] ), .QN(n746) );
  DFFRX1 \CACHE_reg[1][18]  ( .D(n1985), .CK(clk), .RN(n3748), .Q(
        \CACHE[1][18] ), .QN(n745) );
  DFFRX1 \CACHE_reg[1][17]  ( .D(n1984), .CK(clk), .RN(n3748), .Q(
        \CACHE[1][17] ), .QN(n744) );
  DFFRX1 \CACHE_reg[1][16]  ( .D(n1983), .CK(clk), .RN(n3748), .Q(
        \CACHE[1][16] ), .QN(n743) );
  DFFRX1 \CACHE_reg[1][15]  ( .D(n1982), .CK(clk), .RN(n3748), .Q(
        \CACHE[1][15] ), .QN(n742) );
  DFFRX1 \CACHE_reg[1][14]  ( .D(n1981), .CK(clk), .RN(n3748), .Q(
        \CACHE[1][14] ), .QN(n741) );
  DFFRX1 \CACHE_reg[1][13]  ( .D(n1980), .CK(clk), .RN(n3748), .Q(
        \CACHE[1][13] ), .QN(n740) );
  DFFRX1 \CACHE_reg[1][12]  ( .D(n1979), .CK(clk), .RN(n3747), .Q(
        \CACHE[1][12] ), .QN(n739) );
  DFFRX1 \CACHE_reg[1][11]  ( .D(n1978), .CK(clk), .RN(n3747), .Q(
        \CACHE[1][11] ), .QN(n738) );
  DFFRX1 \CACHE_reg[1][10]  ( .D(n1977), .CK(clk), .RN(n3747), .Q(
        \CACHE[1][10] ), .QN(n737) );
  DFFRX1 \CACHE_reg[1][9]  ( .D(n1976), .CK(clk), .RN(n3747), .Q(\CACHE[1][9] ), .QN(n736) );
  DFFRX1 \CACHE_reg[1][8]  ( .D(n1975), .CK(clk), .RN(n3747), .Q(\CACHE[1][8] ), .QN(n735) );
  DFFRX1 \CACHE_reg[1][7]  ( .D(n1974), .CK(clk), .RN(n3747), .Q(\CACHE[1][7] ), .QN(n734) );
  DFFRX1 \CACHE_reg[1][6]  ( .D(n1973), .CK(clk), .RN(n3747), .Q(\CACHE[1][6] ), .QN(n733) );
  DFFRX1 \CACHE_reg[1][5]  ( .D(n1972), .CK(clk), .RN(n3747), .Q(\CACHE[1][5] ), .QN(n732) );
  DFFRX1 \CACHE_reg[1][4]  ( .D(n1971), .CK(clk), .RN(n3747), .Q(\CACHE[1][4] ), .QN(n731) );
  DFFRX1 \CACHE_reg[1][3]  ( .D(n1970), .CK(clk), .RN(n3747), .Q(\CACHE[1][3] ), .QN(n730) );
  DFFRX1 \CACHE_reg[1][2]  ( .D(n1969), .CK(clk), .RN(n3747), .Q(\CACHE[1][2] ), .QN(n729) );
  DFFRX1 \CACHE_reg[1][1]  ( .D(n1968), .CK(clk), .RN(n3747), .Q(\CACHE[1][1] ), .QN(n728) );
  DFFRX1 \CACHE_reg[1][0]  ( .D(n1967), .CK(clk), .RN(n3746), .Q(\CACHE[1][0] ), .QN(n727) );
  DFFRX1 \CACHE_reg[4][118]  ( .D(n2550), .CK(clk), .RN(n3795), .Q(
        \CACHE[4][118] ), .QN(n1310) );
  DFFRX1 \CACHE_reg[4][117]  ( .D(n2549), .CK(clk), .RN(n3795), .Q(
        \CACHE[4][117] ), .QN(n1309) );
  DFFRX1 \CACHE_reg[4][116]  ( .D(n2548), .CK(clk), .RN(n3795), .Q(
        \CACHE[4][116] ), .QN(n1308) );
  DFFRX1 \CACHE_reg[4][115]  ( .D(n2547), .CK(clk), .RN(n3795), .Q(
        \CACHE[4][115] ), .QN(n1307) );
  DFFRX1 \CACHE_reg[4][114]  ( .D(n2546), .CK(clk), .RN(n3795), .Q(
        \CACHE[4][114] ), .QN(n1306) );
  DFFRX1 \CACHE_reg[4][113]  ( .D(n2545), .CK(clk), .RN(n3795), .Q(
        \CACHE[4][113] ), .QN(n1305) );
  DFFRX1 \CACHE_reg[4][112]  ( .D(n2544), .CK(clk), .RN(n3795), .Q(
        \CACHE[4][112] ), .QN(n1304) );
  DFFRX1 \CACHE_reg[4][111]  ( .D(n2543), .CK(clk), .RN(n3794), .Q(
        \CACHE[4][111] ), .QN(n1303) );
  DFFRX1 \CACHE_reg[4][110]  ( .D(n2542), .CK(clk), .RN(n3794), .Q(
        \CACHE[4][110] ), .QN(n1302) );
  DFFRX1 \CACHE_reg[4][109]  ( .D(n2541), .CK(clk), .RN(n3794), .Q(
        \CACHE[4][109] ), .QN(n1301) );
  DFFRX1 \CACHE_reg[4][108]  ( .D(n2540), .CK(clk), .RN(n3794), .Q(
        \CACHE[4][108] ), .QN(n1300) );
  DFFRX1 \CACHE_reg[4][107]  ( .D(n2539), .CK(clk), .RN(n3794), .Q(
        \CACHE[4][107] ), .QN(n1299) );
  DFFRX1 \CACHE_reg[4][106]  ( .D(n2538), .CK(clk), .RN(n3794), .Q(
        \CACHE[4][106] ), .QN(n1298) );
  DFFRX1 \CACHE_reg[4][105]  ( .D(n2537), .CK(clk), .RN(n3794), .Q(
        \CACHE[4][105] ), .QN(n1297) );
  DFFRX1 \CACHE_reg[4][104]  ( .D(n2536), .CK(clk), .RN(n3794), .Q(
        \CACHE[4][104] ), .QN(n1296) );
  DFFRX1 \CACHE_reg[4][103]  ( .D(n2535), .CK(clk), .RN(n3794), .Q(
        \CACHE[4][103] ), .QN(n1295) );
  DFFRX1 \CACHE_reg[4][102]  ( .D(n2534), .CK(clk), .RN(n3794), .Q(
        \CACHE[4][102] ), .QN(n1294) );
  DFFRX1 \CACHE_reg[4][101]  ( .D(n2533), .CK(clk), .RN(n3794), .Q(
        \CACHE[4][101] ), .QN(n1293) );
  DFFRX1 \CACHE_reg[4][100]  ( .D(n2532), .CK(clk), .RN(n3794), .Q(
        \CACHE[4][100] ), .QN(n1292) );
  DFFRX1 \CACHE_reg[4][99]  ( .D(n2531), .CK(clk), .RN(n3793), .Q(
        \CACHE[4][99] ), .QN(n1291) );
  DFFRX1 \CACHE_reg[4][98]  ( .D(n2530), .CK(clk), .RN(n3793), .Q(
        \CACHE[4][98] ), .QN(n1290) );
  DFFRX1 \CACHE_reg[4][97]  ( .D(n2529), .CK(clk), .RN(n3793), .Q(
        \CACHE[4][97] ), .QN(n1289) );
  DFFRX1 \CACHE_reg[4][96]  ( .D(n2528), .CK(clk), .RN(n3793), .Q(
        \CACHE[4][96] ), .QN(n1288) );
  DFFRX1 \CACHE_reg[4][95]  ( .D(n2527), .CK(clk), .RN(n3793), .Q(
        \CACHE[4][95] ), .QN(n1287) );
  DFFRX1 \CACHE_reg[4][94]  ( .D(n2526), .CK(clk), .RN(n3793), .Q(
        \CACHE[4][94] ), .QN(n1286) );
  DFFRX1 \CACHE_reg[4][93]  ( .D(n2525), .CK(clk), .RN(n3793), .Q(
        \CACHE[4][93] ), .QN(n1285) );
  DFFRX1 \CACHE_reg[4][92]  ( .D(n2524), .CK(clk), .RN(n3793), .Q(
        \CACHE[4][92] ), .QN(n1284) );
  DFFRX1 \CACHE_reg[4][91]  ( .D(n2523), .CK(clk), .RN(n3793), .Q(
        \CACHE[4][91] ), .QN(n1283) );
  DFFRX1 \CACHE_reg[4][90]  ( .D(n2522), .CK(clk), .RN(n3793), .Q(
        \CACHE[4][90] ), .QN(n1282) );
  DFFRX1 \CACHE_reg[4][89]  ( .D(n2521), .CK(clk), .RN(n3793), .Q(
        \CACHE[4][89] ), .QN(n1281) );
  DFFRX1 \CACHE_reg[4][88]  ( .D(n2520), .CK(clk), .RN(n3793), .Q(
        \CACHE[4][88] ), .QN(n1280) );
  DFFRX1 \CACHE_reg[4][87]  ( .D(n2519), .CK(clk), .RN(n3792), .Q(
        \CACHE[4][87] ), .QN(n1279) );
  DFFRX1 \CACHE_reg[4][86]  ( .D(n2518), .CK(clk), .RN(n3792), .Q(
        \CACHE[4][86] ), .QN(n1278) );
  DFFRX1 \CACHE_reg[4][85]  ( .D(n2517), .CK(clk), .RN(n3792), .Q(
        \CACHE[4][85] ), .QN(n1277) );
  DFFRX1 \CACHE_reg[4][84]  ( .D(n2516), .CK(clk), .RN(n3792), .Q(
        \CACHE[4][84] ), .QN(n1276) );
  DFFRX1 \CACHE_reg[4][83]  ( .D(n2515), .CK(clk), .RN(n3792), .Q(
        \CACHE[4][83] ), .QN(n1275) );
  DFFRX1 \CACHE_reg[4][82]  ( .D(n2514), .CK(clk), .RN(n3792), .Q(
        \CACHE[4][82] ), .QN(n1274) );
  DFFRX1 \CACHE_reg[4][81]  ( .D(n2513), .CK(clk), .RN(n3792), .Q(
        \CACHE[4][81] ), .QN(n1273) );
  DFFRX1 \CACHE_reg[4][80]  ( .D(n2512), .CK(clk), .RN(n3792), .Q(
        \CACHE[4][80] ), .QN(n1272) );
  DFFRX1 \CACHE_reg[4][79]  ( .D(n2511), .CK(clk), .RN(n3792), .Q(
        \CACHE[4][79] ), .QN(n1271) );
  DFFRX1 \CACHE_reg[4][78]  ( .D(n2510), .CK(clk), .RN(n3792), .Q(
        \CACHE[4][78] ), .QN(n1270) );
  DFFRX1 \CACHE_reg[4][77]  ( .D(n2509), .CK(clk), .RN(n3792), .Q(
        \CACHE[4][77] ), .QN(n1269) );
  DFFRX1 \CACHE_reg[4][76]  ( .D(n2508), .CK(clk), .RN(n3792), .Q(
        \CACHE[4][76] ), .QN(n1268) );
  DFFRX1 \CACHE_reg[4][75]  ( .D(n2507), .CK(clk), .RN(n3791), .Q(
        \CACHE[4][75] ), .QN(n1267) );
  DFFRX1 \CACHE_reg[4][74]  ( .D(n2506), .CK(clk), .RN(n3791), .Q(
        \CACHE[4][74] ), .QN(n1266) );
  DFFRX1 \CACHE_reg[4][73]  ( .D(n2505), .CK(clk), .RN(n3791), .Q(
        \CACHE[4][73] ), .QN(n1265) );
  DFFRX1 \CACHE_reg[4][72]  ( .D(n2504), .CK(clk), .RN(n3791), .Q(
        \CACHE[4][72] ), .QN(n1264) );
  DFFRX1 \CACHE_reg[4][71]  ( .D(n2503), .CK(clk), .RN(n3791), .Q(
        \CACHE[4][71] ), .QN(n1263) );
  DFFRX1 \CACHE_reg[4][70]  ( .D(n2502), .CK(clk), .RN(n3791), .Q(
        \CACHE[4][70] ), .QN(n1262) );
  DFFRX1 \CACHE_reg[4][69]  ( .D(n2501), .CK(clk), .RN(n3791), .Q(
        \CACHE[4][69] ), .QN(n1261) );
  DFFRX1 \CACHE_reg[4][68]  ( .D(n2500), .CK(clk), .RN(n3791), .Q(
        \CACHE[4][68] ), .QN(n1260) );
  DFFRX1 \CACHE_reg[4][67]  ( .D(n2499), .CK(clk), .RN(n3791), .Q(
        \CACHE[4][67] ), .QN(n1259) );
  DFFRX1 \CACHE_reg[4][66]  ( .D(n2498), .CK(clk), .RN(n3791), .Q(
        \CACHE[4][66] ), .QN(n1258) );
  DFFRX1 \CACHE_reg[4][65]  ( .D(n2497), .CK(clk), .RN(n3791), .Q(
        \CACHE[4][65] ), .QN(n1257) );
  DFFRX1 \CACHE_reg[4][64]  ( .D(n2496), .CK(clk), .RN(n3791), .Q(
        \CACHE[4][64] ), .QN(n1256) );
  DFFRX1 \CACHE_reg[4][63]  ( .D(n2495), .CK(clk), .RN(n3790), .Q(
        \CACHE[4][63] ), .QN(n1255) );
  DFFRX1 \CACHE_reg[4][62]  ( .D(n2494), .CK(clk), .RN(n3790), .Q(
        \CACHE[4][62] ), .QN(n1254) );
  DFFRX1 \CACHE_reg[4][61]  ( .D(n2493), .CK(clk), .RN(n3790), .Q(
        \CACHE[4][61] ), .QN(n1253) );
  DFFRX1 \CACHE_reg[4][60]  ( .D(n2492), .CK(clk), .RN(n3790), .Q(
        \CACHE[4][60] ), .QN(n1252) );
  DFFRX1 \CACHE_reg[4][59]  ( .D(n2491), .CK(clk), .RN(n3790), .Q(
        \CACHE[4][59] ), .QN(n1251) );
  DFFRX1 \CACHE_reg[4][58]  ( .D(n2490), .CK(clk), .RN(n3790), .Q(
        \CACHE[4][58] ), .QN(n1250) );
  DFFRX1 \CACHE_reg[4][57]  ( .D(n2489), .CK(clk), .RN(n3790), .Q(
        \CACHE[4][57] ), .QN(n1249) );
  DFFRX1 \CACHE_reg[4][56]  ( .D(n2488), .CK(clk), .RN(n3790), .Q(
        \CACHE[4][56] ), .QN(n1248) );
  DFFRX1 \CACHE_reg[4][55]  ( .D(n2487), .CK(clk), .RN(n3790), .Q(
        \CACHE[4][55] ), .QN(n1247) );
  DFFRX1 \CACHE_reg[4][54]  ( .D(n2486), .CK(clk), .RN(n3790), .Q(
        \CACHE[4][54] ), .QN(n1246) );
  DFFRX1 \CACHE_reg[4][53]  ( .D(n2485), .CK(clk), .RN(n3790), .Q(
        \CACHE[4][53] ), .QN(n1245) );
  DFFRX1 \CACHE_reg[4][52]  ( .D(n2484), .CK(clk), .RN(n3790), .Q(
        \CACHE[4][52] ), .QN(n1244) );
  DFFRX1 \CACHE_reg[4][51]  ( .D(n2483), .CK(clk), .RN(n3789), .Q(
        \CACHE[4][51] ), .QN(n1243) );
  DFFRX1 \CACHE_reg[4][50]  ( .D(n2482), .CK(clk), .RN(n3789), .Q(
        \CACHE[4][50] ), .QN(n1242) );
  DFFRX1 \CACHE_reg[4][49]  ( .D(n2481), .CK(clk), .RN(n3789), .Q(
        \CACHE[4][49] ), .QN(n1241) );
  DFFRX1 \CACHE_reg[4][48]  ( .D(n2480), .CK(clk), .RN(n3789), .Q(
        \CACHE[4][48] ), .QN(n1240) );
  DFFRX1 \CACHE_reg[4][47]  ( .D(n2479), .CK(clk), .RN(n3789), .Q(
        \CACHE[4][47] ), .QN(n1239) );
  DFFRX1 \CACHE_reg[4][46]  ( .D(n2478), .CK(clk), .RN(n3789), .Q(
        \CACHE[4][46] ), .QN(n1238) );
  DFFRX1 \CACHE_reg[4][45]  ( .D(n2477), .CK(clk), .RN(n3789), .Q(
        \CACHE[4][45] ), .QN(n1237) );
  DFFRX1 \CACHE_reg[4][44]  ( .D(n2476), .CK(clk), .RN(n3789), .Q(
        \CACHE[4][44] ), .QN(n1236) );
  DFFRX1 \CACHE_reg[4][43]  ( .D(n2475), .CK(clk), .RN(n3789), .Q(
        \CACHE[4][43] ), .QN(n1235) );
  DFFRX1 \CACHE_reg[4][42]  ( .D(n2474), .CK(clk), .RN(n3789), .Q(
        \CACHE[4][42] ), .QN(n1234) );
  DFFRX1 \CACHE_reg[4][41]  ( .D(n2473), .CK(clk), .RN(n3789), .Q(
        \CACHE[4][41] ), .QN(n1233) );
  DFFRX1 \CACHE_reg[4][40]  ( .D(n2472), .CK(clk), .RN(n3789), .Q(
        \CACHE[4][40] ), .QN(n1232) );
  DFFRX1 \CACHE_reg[4][39]  ( .D(n2471), .CK(clk), .RN(n3788), .Q(
        \CACHE[4][39] ), .QN(n1231) );
  DFFRX1 \CACHE_reg[4][38]  ( .D(n2470), .CK(clk), .RN(n3788), .Q(
        \CACHE[4][38] ), .QN(n1230) );
  DFFRX1 \CACHE_reg[4][37]  ( .D(n2469), .CK(clk), .RN(n3788), .Q(
        \CACHE[4][37] ), .QN(n1229) );
  DFFRX1 \CACHE_reg[4][36]  ( .D(n2468), .CK(clk), .RN(n3788), .Q(
        \CACHE[4][36] ), .QN(n1228) );
  DFFRX1 \CACHE_reg[4][35]  ( .D(n2467), .CK(clk), .RN(n3788), .Q(
        \CACHE[4][35] ), .QN(n1227) );
  DFFRX1 \CACHE_reg[4][34]  ( .D(n2466), .CK(clk), .RN(n3788), .Q(
        \CACHE[4][34] ), .QN(n1226) );
  DFFRX1 \CACHE_reg[4][33]  ( .D(n2465), .CK(clk), .RN(n3788), .Q(
        \CACHE[4][33] ), .QN(n1225) );
  DFFRX1 \CACHE_reg[4][32]  ( .D(n2464), .CK(clk), .RN(n3788), .Q(
        \CACHE[4][32] ), .QN(n1224) );
  DFFRX1 \CACHE_reg[4][31]  ( .D(n2463), .CK(clk), .RN(n3788), .Q(
        \CACHE[4][31] ), .QN(n1223) );
  DFFRX1 \CACHE_reg[4][30]  ( .D(n2462), .CK(clk), .RN(n3788), .Q(
        \CACHE[4][30] ), .QN(n1222) );
  DFFRX1 \CACHE_reg[4][29]  ( .D(n2461), .CK(clk), .RN(n3788), .Q(
        \CACHE[4][29] ), .QN(n1221) );
  DFFRX1 \CACHE_reg[4][28]  ( .D(n2460), .CK(clk), .RN(n3788), .Q(
        \CACHE[4][28] ), .QN(n1220) );
  DFFRX1 \CACHE_reg[4][27]  ( .D(n2459), .CK(clk), .RN(n3787), .Q(
        \CACHE[4][27] ), .QN(n1219) );
  DFFRX1 \CACHE_reg[4][26]  ( .D(n2458), .CK(clk), .RN(n3787), .Q(
        \CACHE[4][26] ), .QN(n1218) );
  DFFRX1 \CACHE_reg[4][25]  ( .D(n2457), .CK(clk), .RN(n3787), .Q(
        \CACHE[4][25] ), .QN(n1217) );
  DFFRX1 \CACHE_reg[4][24]  ( .D(n2456), .CK(clk), .RN(n3787), .Q(
        \CACHE[4][24] ), .QN(n1216) );
  DFFRX1 \CACHE_reg[4][23]  ( .D(n2455), .CK(clk), .RN(n3787), .Q(
        \CACHE[4][23] ), .QN(n1215) );
  DFFRX1 \CACHE_reg[4][22]  ( .D(n2454), .CK(clk), .RN(n3787), .Q(
        \CACHE[4][22] ), .QN(n1214) );
  DFFRX1 \CACHE_reg[4][21]  ( .D(n2453), .CK(clk), .RN(n3787), .Q(
        \CACHE[4][21] ), .QN(n1213) );
  DFFRX1 \CACHE_reg[4][20]  ( .D(n2452), .CK(clk), .RN(n3787), .Q(
        \CACHE[4][20] ), .QN(n1212) );
  DFFRX1 \CACHE_reg[4][19]  ( .D(n2451), .CK(clk), .RN(n3787), .Q(
        \CACHE[4][19] ), .QN(n1211) );
  DFFRX1 \CACHE_reg[4][18]  ( .D(n2450), .CK(clk), .RN(n3787), .Q(
        \CACHE[4][18] ), .QN(n1210) );
  DFFRX1 \CACHE_reg[4][17]  ( .D(n2449), .CK(clk), .RN(n3787), .Q(
        \CACHE[4][17] ), .QN(n1209) );
  DFFRX1 \CACHE_reg[4][16]  ( .D(n2448), .CK(clk), .RN(n3787), .Q(
        \CACHE[4][16] ), .QN(n1208) );
  DFFRX1 \CACHE_reg[4][15]  ( .D(n2447), .CK(clk), .RN(n3786), .Q(
        \CACHE[4][15] ), .QN(n1207) );
  DFFRX1 \CACHE_reg[4][14]  ( .D(n2446), .CK(clk), .RN(n3786), .Q(
        \CACHE[4][14] ), .QN(n1206) );
  DFFRX1 \CACHE_reg[4][13]  ( .D(n2445), .CK(clk), .RN(n3786), .Q(
        \CACHE[4][13] ), .QN(n1205) );
  DFFRX1 \CACHE_reg[4][12]  ( .D(n2444), .CK(clk), .RN(n3786), .Q(
        \CACHE[4][12] ), .QN(n1204) );
  DFFRX1 \CACHE_reg[4][11]  ( .D(n2443), .CK(clk), .RN(n3786), .Q(
        \CACHE[4][11] ), .QN(n1203) );
  DFFRX1 \CACHE_reg[4][10]  ( .D(n2442), .CK(clk), .RN(n3786), .Q(
        \CACHE[4][10] ), .QN(n1202) );
  DFFRX1 \CACHE_reg[4][9]  ( .D(n2441), .CK(clk), .RN(n3786), .Q(\CACHE[4][9] ), .QN(n1201) );
  DFFRX1 \CACHE_reg[4][8]  ( .D(n2440), .CK(clk), .RN(n3786), .Q(\CACHE[4][8] ), .QN(n1200) );
  DFFRX1 \CACHE_reg[4][7]  ( .D(n2439), .CK(clk), .RN(n3786), .Q(\CACHE[4][7] ), .QN(n1199) );
  DFFRX1 \CACHE_reg[4][6]  ( .D(n2438), .CK(clk), .RN(n3786), .Q(\CACHE[4][6] ), .QN(n1198) );
  DFFRX1 \CACHE_reg[4][5]  ( .D(n2437), .CK(clk), .RN(n3786), .Q(\CACHE[4][5] ), .QN(n1197) );
  DFFRX1 \CACHE_reg[4][4]  ( .D(n2436), .CK(clk), .RN(n3786), .Q(\CACHE[4][4] ), .QN(n1196) );
  DFFRX1 \CACHE_reg[4][3]  ( .D(n2435), .CK(clk), .RN(n3785), .Q(\CACHE[4][3] ), .QN(n1195) );
  DFFRX1 \CACHE_reg[4][2]  ( .D(n2434), .CK(clk), .RN(n3785), .Q(\CACHE[4][2] ), .QN(n1194) );
  DFFRX1 \CACHE_reg[4][1]  ( .D(n2433), .CK(clk), .RN(n3785), .Q(\CACHE[4][1] ), .QN(n1193) );
  DFFRX1 \CACHE_reg[4][0]  ( .D(n2432), .CK(clk), .RN(n3785), .Q(\CACHE[4][0] ), .QN(n1192) );
  DFFRX1 \CACHE_reg[0][118]  ( .D(n1930), .CK(clk), .RN(n3743), .Q(
        \CACHE[0][118] ), .QN(n690) );
  DFFRX1 \CACHE_reg[0][117]  ( .D(n1929), .CK(clk), .RN(n3743), .Q(
        \CACHE[0][117] ), .QN(n689) );
  DFFRX1 \CACHE_reg[0][116]  ( .D(n1928), .CK(clk), .RN(n3743), .Q(
        \CACHE[0][116] ), .QN(n688) );
  DFFRX1 \CACHE_reg[0][115]  ( .D(n1927), .CK(clk), .RN(n3743), .Q(
        \CACHE[0][115] ), .QN(n687) );
  DFFRX1 \CACHE_reg[0][114]  ( .D(n1926), .CK(clk), .RN(n3743), .Q(
        \CACHE[0][114] ), .QN(n686) );
  DFFRX1 \CACHE_reg[0][113]  ( .D(n1925), .CK(clk), .RN(n3743), .Q(
        \CACHE[0][113] ), .QN(n685) );
  DFFRX1 \CACHE_reg[0][112]  ( .D(n1924), .CK(clk), .RN(n3743), .Q(
        \CACHE[0][112] ), .QN(n684) );
  DFFRX1 \CACHE_reg[0][111]  ( .D(n1923), .CK(clk), .RN(n3743), .Q(
        \CACHE[0][111] ), .QN(n683) );
  DFFRX1 \CACHE_reg[0][110]  ( .D(n1922), .CK(clk), .RN(n3743), .Q(
        \CACHE[0][110] ), .QN(n682) );
  DFFRX1 \CACHE_reg[0][109]  ( .D(n1921), .CK(clk), .RN(n3743), .Q(
        \CACHE[0][109] ), .QN(n681) );
  DFFRX1 \CACHE_reg[0][108]  ( .D(n1920), .CK(clk), .RN(n3743), .Q(
        \CACHE[0][108] ), .QN(n680) );
  DFFRX1 \CACHE_reg[0][107]  ( .D(n1919), .CK(clk), .RN(n3742), .Q(
        \CACHE[0][107] ), .QN(n679) );
  DFFRX1 \CACHE_reg[0][106]  ( .D(n1918), .CK(clk), .RN(n3742), .Q(
        \CACHE[0][106] ), .QN(n678) );
  DFFRX1 \CACHE_reg[0][105]  ( .D(n1917), .CK(clk), .RN(n3742), .Q(
        \CACHE[0][105] ), .QN(n677) );
  DFFRX1 \CACHE_reg[0][104]  ( .D(n1916), .CK(clk), .RN(n3742), .Q(
        \CACHE[0][104] ), .QN(n676) );
  DFFRX1 \CACHE_reg[0][103]  ( .D(n1915), .CK(clk), .RN(n3742), .Q(
        \CACHE[0][103] ), .QN(n675) );
  DFFRX1 \CACHE_reg[0][102]  ( .D(n1914), .CK(clk), .RN(n3742), .Q(
        \CACHE[0][102] ), .QN(n674) );
  DFFRX1 \CACHE_reg[0][101]  ( .D(n1913), .CK(clk), .RN(n3742), .Q(
        \CACHE[0][101] ), .QN(n673) );
  DFFRX1 \CACHE_reg[0][100]  ( .D(n1912), .CK(clk), .RN(n3742), .Q(
        \CACHE[0][100] ), .QN(n672) );
  DFFRX1 \CACHE_reg[0][99]  ( .D(n1911), .CK(clk), .RN(n3742), .Q(
        \CACHE[0][99] ), .QN(n671) );
  DFFRX1 \CACHE_reg[0][98]  ( .D(n1910), .CK(clk), .RN(n3742), .Q(
        \CACHE[0][98] ), .QN(n670) );
  DFFRX1 \CACHE_reg[0][97]  ( .D(n1909), .CK(clk), .RN(n3742), .Q(
        \CACHE[0][97] ), .QN(n669) );
  DFFRX1 \CACHE_reg[0][96]  ( .D(n1908), .CK(clk), .RN(n3742), .Q(
        \CACHE[0][96] ), .QN(n668) );
  DFFRX1 \CACHE_reg[0][95]  ( .D(n1907), .CK(clk), .RN(n3741), .Q(
        \CACHE[0][95] ), .QN(n667) );
  DFFRX1 \CACHE_reg[0][94]  ( .D(n1906), .CK(clk), .RN(n3741), .Q(
        \CACHE[0][94] ), .QN(n666) );
  DFFRX1 \CACHE_reg[0][93]  ( .D(n1905), .CK(clk), .RN(n3741), .Q(
        \CACHE[0][93] ), .QN(n665) );
  DFFRX1 \CACHE_reg[0][92]  ( .D(n1904), .CK(clk), .RN(n3741), .Q(
        \CACHE[0][92] ), .QN(n664) );
  DFFRX1 \CACHE_reg[0][91]  ( .D(n1903), .CK(clk), .RN(n3741), .Q(
        \CACHE[0][91] ), .QN(n663) );
  DFFRX1 \CACHE_reg[0][90]  ( .D(n1902), .CK(clk), .RN(n3741), .Q(
        \CACHE[0][90] ), .QN(n662) );
  DFFRX1 \CACHE_reg[0][89]  ( .D(n1901), .CK(clk), .RN(n3741), .Q(
        \CACHE[0][89] ), .QN(n661) );
  DFFRX1 \CACHE_reg[0][88]  ( .D(n1900), .CK(clk), .RN(n3741), .Q(
        \CACHE[0][88] ), .QN(n660) );
  DFFRX1 \CACHE_reg[0][87]  ( .D(n1899), .CK(clk), .RN(n3741), .Q(
        \CACHE[0][87] ), .QN(n659) );
  DFFRX1 \CACHE_reg[0][86]  ( .D(n1898), .CK(clk), .RN(n3741), .Q(
        \CACHE[0][86] ), .QN(n658) );
  DFFRX1 \CACHE_reg[0][85]  ( .D(n1897), .CK(clk), .RN(n3741), .Q(
        \CACHE[0][85] ), .QN(n657) );
  DFFRX1 \CACHE_reg[0][84]  ( .D(n1896), .CK(clk), .RN(n3741), .Q(
        \CACHE[0][84] ), .QN(n656) );
  DFFRX1 \CACHE_reg[0][83]  ( .D(n1895), .CK(clk), .RN(n3740), .Q(
        \CACHE[0][83] ), .QN(n655) );
  DFFRX1 \CACHE_reg[0][82]  ( .D(n1894), .CK(clk), .RN(n3740), .Q(
        \CACHE[0][82] ), .QN(n654) );
  DFFRX1 \CACHE_reg[0][81]  ( .D(n1893), .CK(clk), .RN(n3740), .Q(
        \CACHE[0][81] ), .QN(n653) );
  DFFRX1 \CACHE_reg[0][80]  ( .D(n1892), .CK(clk), .RN(n3740), .Q(
        \CACHE[0][80] ), .QN(n652) );
  DFFRX1 \CACHE_reg[0][79]  ( .D(n1891), .CK(clk), .RN(n3740), .Q(
        \CACHE[0][79] ), .QN(n651) );
  DFFRX1 \CACHE_reg[0][78]  ( .D(n1890), .CK(clk), .RN(n3740), .Q(
        \CACHE[0][78] ), .QN(n650) );
  DFFRX1 \CACHE_reg[0][77]  ( .D(n1889), .CK(clk), .RN(n3740), .Q(
        \CACHE[0][77] ), .QN(n649) );
  DFFRX1 \CACHE_reg[0][76]  ( .D(n1888), .CK(clk), .RN(n3740), .Q(
        \CACHE[0][76] ), .QN(n648) );
  DFFRX1 \CACHE_reg[0][75]  ( .D(n1887), .CK(clk), .RN(n3740), .Q(
        \CACHE[0][75] ), .QN(n647) );
  DFFRX1 \CACHE_reg[0][74]  ( .D(n1886), .CK(clk), .RN(n3740), .Q(
        \CACHE[0][74] ), .QN(n646) );
  DFFRX1 \CACHE_reg[0][73]  ( .D(n1885), .CK(clk), .RN(n3740), .Q(
        \CACHE[0][73] ), .QN(n645) );
  DFFRX1 \CACHE_reg[0][72]  ( .D(n1884), .CK(clk), .RN(n3740), .Q(
        \CACHE[0][72] ), .QN(n644) );
  DFFRX1 \CACHE_reg[0][71]  ( .D(n1883), .CK(clk), .RN(n3739), .Q(
        \CACHE[0][71] ), .QN(n643) );
  DFFRX1 \CACHE_reg[0][70]  ( .D(n1882), .CK(clk), .RN(n3739), .Q(
        \CACHE[0][70] ), .QN(n642) );
  DFFRX1 \CACHE_reg[0][69]  ( .D(n1881), .CK(clk), .RN(n3739), .Q(
        \CACHE[0][69] ), .QN(n641) );
  DFFRX1 \CACHE_reg[0][68]  ( .D(n1880), .CK(clk), .RN(n3739), .Q(
        \CACHE[0][68] ), .QN(n640) );
  DFFRX1 \CACHE_reg[0][67]  ( .D(n1879), .CK(clk), .RN(n3739), .Q(
        \CACHE[0][67] ), .QN(n639) );
  DFFRX1 \CACHE_reg[0][66]  ( .D(n1878), .CK(clk), .RN(n3739), .Q(
        \CACHE[0][66] ), .QN(n638) );
  DFFRX1 \CACHE_reg[0][65]  ( .D(n1877), .CK(clk), .RN(n3739), .Q(
        \CACHE[0][65] ), .QN(n637) );
  DFFRX1 \CACHE_reg[0][64]  ( .D(n1876), .CK(clk), .RN(n3739), .Q(
        \CACHE[0][64] ), .QN(n636) );
  DFFRX1 \CACHE_reg[0][63]  ( .D(n1875), .CK(clk), .RN(n3739), .Q(
        \CACHE[0][63] ), .QN(n635) );
  DFFRX1 \CACHE_reg[0][62]  ( .D(n1874), .CK(clk), .RN(n3739), .Q(
        \CACHE[0][62] ), .QN(n634) );
  DFFRX1 \CACHE_reg[0][61]  ( .D(n1873), .CK(clk), .RN(n3739), .Q(
        \CACHE[0][61] ), .QN(n633) );
  DFFRX1 \CACHE_reg[0][60]  ( .D(n1872), .CK(clk), .RN(n3739), .Q(
        \CACHE[0][60] ), .QN(n632) );
  DFFRX1 \CACHE_reg[0][59]  ( .D(n1871), .CK(clk), .RN(n3738), .Q(
        \CACHE[0][59] ), .QN(n631) );
  DFFRX1 \CACHE_reg[0][58]  ( .D(n1870), .CK(clk), .RN(n3738), .Q(
        \CACHE[0][58] ), .QN(n630) );
  DFFRX1 \CACHE_reg[0][57]  ( .D(n1869), .CK(clk), .RN(n3738), .Q(
        \CACHE[0][57] ), .QN(n629) );
  DFFRX1 \CACHE_reg[0][56]  ( .D(n1868), .CK(clk), .RN(n3738), .Q(
        \CACHE[0][56] ), .QN(n628) );
  DFFRX1 \CACHE_reg[0][55]  ( .D(n1867), .CK(clk), .RN(n3738), .Q(
        \CACHE[0][55] ), .QN(n627) );
  DFFRX1 \CACHE_reg[0][54]  ( .D(n1866), .CK(clk), .RN(n3738), .Q(
        \CACHE[0][54] ), .QN(n626) );
  DFFRX1 \CACHE_reg[0][53]  ( .D(n1865), .CK(clk), .RN(n3738), .Q(
        \CACHE[0][53] ), .QN(n625) );
  DFFRX1 \CACHE_reg[0][52]  ( .D(n1864), .CK(clk), .RN(n3738), .Q(
        \CACHE[0][52] ), .QN(n624) );
  DFFRX1 \CACHE_reg[0][51]  ( .D(n1863), .CK(clk), .RN(n3738), .Q(
        \CACHE[0][51] ), .QN(n623) );
  DFFRX1 \CACHE_reg[0][50]  ( .D(n1862), .CK(clk), .RN(n3738), .Q(
        \CACHE[0][50] ), .QN(n622) );
  DFFRX1 \CACHE_reg[0][49]  ( .D(n1861), .CK(clk), .RN(n3738), .Q(
        \CACHE[0][49] ), .QN(n621) );
  DFFRX1 \CACHE_reg[0][48]  ( .D(n1860), .CK(clk), .RN(n3738), .Q(
        \CACHE[0][48] ), .QN(n620) );
  DFFRX1 \CACHE_reg[0][47]  ( .D(n1859), .CK(clk), .RN(n3737), .Q(
        \CACHE[0][47] ), .QN(n619) );
  DFFRX1 \CACHE_reg[0][46]  ( .D(n1858), .CK(clk), .RN(n3737), .Q(
        \CACHE[0][46] ), .QN(n618) );
  DFFRX1 \CACHE_reg[0][45]  ( .D(n1857), .CK(clk), .RN(n3737), .Q(
        \CACHE[0][45] ), .QN(n617) );
  DFFRX1 \CACHE_reg[0][44]  ( .D(n1856), .CK(clk), .RN(n3737), .Q(
        \CACHE[0][44] ), .QN(n616) );
  DFFRX1 \CACHE_reg[0][43]  ( .D(n1855), .CK(clk), .RN(n3737), .Q(
        \CACHE[0][43] ), .QN(n615) );
  DFFRX1 \CACHE_reg[0][42]  ( .D(n1854), .CK(clk), .RN(n3737), .Q(
        \CACHE[0][42] ), .QN(n614) );
  DFFRX1 \CACHE_reg[0][41]  ( .D(n1853), .CK(clk), .RN(n3737), .Q(
        \CACHE[0][41] ), .QN(n613) );
  DFFRX1 \CACHE_reg[0][40]  ( .D(n1852), .CK(clk), .RN(n3737), .Q(
        \CACHE[0][40] ), .QN(n612) );
  DFFRX1 \CACHE_reg[0][39]  ( .D(n1851), .CK(clk), .RN(n3737), .Q(
        \CACHE[0][39] ), .QN(n611) );
  DFFRX1 \CACHE_reg[0][38]  ( .D(n1850), .CK(clk), .RN(n3737), .Q(
        \CACHE[0][38] ), .QN(n610) );
  DFFRX1 \CACHE_reg[0][37]  ( .D(n1849), .CK(clk), .RN(n3737), .Q(
        \CACHE[0][37] ), .QN(n609) );
  DFFRX1 \CACHE_reg[0][35]  ( .D(n1847), .CK(clk), .RN(n3736), .Q(
        \CACHE[0][35] ), .QN(n607) );
  DFFRX1 \CACHE_reg[0][34]  ( .D(n1846), .CK(clk), .RN(n3736), .Q(
        \CACHE[0][34] ), .QN(n606) );
  DFFRX1 \CACHE_reg[0][33]  ( .D(n1845), .CK(clk), .RN(n3736), .Q(
        \CACHE[0][33] ), .QN(n605) );
  DFFRX1 \CACHE_reg[0][31]  ( .D(n1843), .CK(clk), .RN(n3736), .Q(
        \CACHE[0][31] ), .QN(n603) );
  DFFRX1 \CACHE_reg[0][30]  ( .D(n1842), .CK(clk), .RN(n3736), .Q(
        \CACHE[0][30] ), .QN(n602) );
  DFFRX1 \CACHE_reg[0][29]  ( .D(n1841), .CK(clk), .RN(n3736), .Q(
        \CACHE[0][29] ), .QN(n601) );
  DFFRX1 \CACHE_reg[0][28]  ( .D(n1840), .CK(clk), .RN(n3736), .Q(
        \CACHE[0][28] ), .QN(n600) );
  DFFRX1 \CACHE_reg[0][27]  ( .D(n1839), .CK(clk), .RN(n3736), .Q(
        \CACHE[0][27] ), .QN(n599) );
  DFFRX1 \CACHE_reg[0][26]  ( .D(n1838), .CK(clk), .RN(n3736), .Q(
        \CACHE[0][26] ), .QN(n598) );
  DFFRX1 \CACHE_reg[0][25]  ( .D(n1837), .CK(clk), .RN(n3736), .Q(
        \CACHE[0][25] ), .QN(n597) );
  DFFRX1 \CACHE_reg[0][24]  ( .D(n1836), .CK(clk), .RN(n3736), .Q(
        \CACHE[0][24] ), .QN(n596) );
  DFFRX1 \CACHE_reg[0][23]  ( .D(n1835), .CK(clk), .RN(n3735), .Q(
        \CACHE[0][23] ), .QN(n595) );
  DFFRX1 \CACHE_reg[0][22]  ( .D(n1834), .CK(clk), .RN(n3735), .Q(
        \CACHE[0][22] ), .QN(n594) );
  DFFRX1 \CACHE_reg[0][21]  ( .D(n1833), .CK(clk), .RN(n3735), .Q(
        \CACHE[0][21] ), .QN(n593) );
  DFFRX1 \CACHE_reg[0][20]  ( .D(n1832), .CK(clk), .RN(n3735), .Q(
        \CACHE[0][20] ), .QN(n592) );
  DFFRX1 \CACHE_reg[0][19]  ( .D(n1831), .CK(clk), .RN(n3735), .Q(
        \CACHE[0][19] ), .QN(n591) );
  DFFRX1 \CACHE_reg[0][18]  ( .D(n1830), .CK(clk), .RN(n3735), .Q(
        \CACHE[0][18] ), .QN(n590) );
  DFFRX1 \CACHE_reg[0][17]  ( .D(n1829), .CK(clk), .RN(n3735), .Q(
        \CACHE[0][17] ), .QN(n589) );
  DFFRX1 \CACHE_reg[0][16]  ( .D(n1828), .CK(clk), .RN(n3735), .Q(
        \CACHE[0][16] ), .QN(n588) );
  DFFRX1 \CACHE_reg[0][15]  ( .D(n1827), .CK(clk), .RN(n3735), .Q(
        \CACHE[0][15] ), .QN(n587) );
  DFFRX1 \CACHE_reg[0][14]  ( .D(n1826), .CK(clk), .RN(n3735), .Q(
        \CACHE[0][14] ), .QN(n586) );
  DFFRX1 \CACHE_reg[0][13]  ( .D(n1825), .CK(clk), .RN(n3735), .Q(
        \CACHE[0][13] ), .QN(n585) );
  DFFRX1 \CACHE_reg[0][12]  ( .D(n1824), .CK(clk), .RN(n3735), .Q(
        \CACHE[0][12] ), .QN(n584) );
  DFFRX1 \CACHE_reg[0][11]  ( .D(n1823), .CK(clk), .RN(n3734), .Q(
        \CACHE[0][11] ), .QN(n583) );
  DFFRX1 \CACHE_reg[0][10]  ( .D(n1822), .CK(clk), .RN(n3734), .Q(
        \CACHE[0][10] ), .QN(n582) );
  DFFRX1 \CACHE_reg[0][9]  ( .D(n1821), .CK(clk), .RN(n3734), .Q(\CACHE[0][9] ), .QN(n581) );
  DFFRX1 \CACHE_reg[0][8]  ( .D(n1820), .CK(clk), .RN(n3734), .Q(\CACHE[0][8] ), .QN(n580) );
  DFFRX1 \CACHE_reg[0][7]  ( .D(n1819), .CK(clk), .RN(n3734), .Q(\CACHE[0][7] ), .QN(n579) );
  DFFRX1 \CACHE_reg[0][6]  ( .D(n1818), .CK(clk), .RN(n3734), .Q(\CACHE[0][6] ), .QN(n578) );
  DFFRX1 \CACHE_reg[0][5]  ( .D(n1817), .CK(clk), .RN(n3734), .Q(\CACHE[0][5] ), .QN(n577) );
  DFFRX1 \CACHE_reg[0][4]  ( .D(n1816), .CK(clk), .RN(n3734), .Q(\CACHE[0][4] ), .QN(n576) );
  DFFRX1 \CACHE_reg[0][3]  ( .D(n1815), .CK(clk), .RN(n3734), .Q(\CACHE[0][3] ), .QN(n575) );
  DFFRX1 \CACHE_reg[0][2]  ( .D(n1814), .CK(clk), .RN(n3734), .Q(\CACHE[0][2] ), .QN(n574) );
  DFFRX1 \CACHE_reg[0][1]  ( .D(n1813), .CK(clk), .RN(n3734), .Q(\CACHE[0][1] ), .QN(n573) );
  DFFRX1 \CACHE_reg[0][0]  ( .D(n1812), .CK(clk), .RN(n3734), .Q(\CACHE[0][0] ), .QN(n572) );
  DFFRX1 \CACHE_reg[6][118]  ( .D(n2860), .CK(clk), .RN(n3821), .Q(
        \CACHE[6][118] ), .QN(n1620) );
  DFFRX1 \CACHE_reg[6][117]  ( .D(n2859), .CK(clk), .RN(n3821), .Q(
        \CACHE[6][117] ), .QN(n1619) );
  DFFRX1 \CACHE_reg[6][116]  ( .D(n2858), .CK(clk), .RN(n3821), .Q(
        \CACHE[6][116] ), .QN(n1618) );
  DFFRX1 \CACHE_reg[6][115]  ( .D(n2857), .CK(clk), .RN(n3821), .Q(
        \CACHE[6][115] ), .QN(n1617) );
  DFFRX1 \CACHE_reg[6][114]  ( .D(n2856), .CK(clk), .RN(n3821), .Q(
        \CACHE[6][114] ), .QN(n1616) );
  DFFRX1 \CACHE_reg[6][113]  ( .D(n2855), .CK(clk), .RN(n3820), .Q(
        \CACHE[6][113] ), .QN(n1615) );
  DFFRX1 \CACHE_reg[6][112]  ( .D(n2854), .CK(clk), .RN(n3820), .Q(
        \CACHE[6][112] ), .QN(n1614) );
  DFFRX1 \CACHE_reg[6][111]  ( .D(n2853), .CK(clk), .RN(n3820), .Q(
        \CACHE[6][111] ), .QN(n1613) );
  DFFRX1 \CACHE_reg[6][110]  ( .D(n2852), .CK(clk), .RN(n3820), .Q(
        \CACHE[6][110] ), .QN(n1612) );
  DFFRX1 \CACHE_reg[6][109]  ( .D(n2851), .CK(clk), .RN(n3820), .Q(
        \CACHE[6][109] ), .QN(n1611) );
  DFFRX1 \CACHE_reg[6][108]  ( .D(n2850), .CK(clk), .RN(n3820), .Q(
        \CACHE[6][108] ), .QN(n1610) );
  DFFRX1 \CACHE_reg[6][107]  ( .D(n2849), .CK(clk), .RN(n3820), .Q(
        \CACHE[6][107] ), .QN(n1609) );
  DFFRX1 \CACHE_reg[6][106]  ( .D(n2848), .CK(clk), .RN(n3820), .Q(
        \CACHE[6][106] ), .QN(n1608) );
  DFFRX1 \CACHE_reg[6][105]  ( .D(n2847), .CK(clk), .RN(n3820), .Q(
        \CACHE[6][105] ), .QN(n1607) );
  DFFRX1 \CACHE_reg[6][104]  ( .D(n2846), .CK(clk), .RN(n3820), .Q(
        \CACHE[6][104] ), .QN(n1606) );
  DFFRX1 \CACHE_reg[6][103]  ( .D(n2845), .CK(clk), .RN(n3820), .Q(
        \CACHE[6][103] ), .QN(n1605) );
  DFFRX1 \CACHE_reg[6][102]  ( .D(n2844), .CK(clk), .RN(n3820), .Q(
        \CACHE[6][102] ), .QN(n1604) );
  DFFRX1 \CACHE_reg[6][101]  ( .D(n2843), .CK(clk), .RN(n3819), .Q(
        \CACHE[6][101] ), .QN(n1603) );
  DFFRX1 \CACHE_reg[6][100]  ( .D(n2842), .CK(clk), .RN(n3819), .Q(
        \CACHE[6][100] ), .QN(n1602) );
  DFFRX1 \CACHE_reg[6][99]  ( .D(n2841), .CK(clk), .RN(n3819), .Q(
        \CACHE[6][99] ), .QN(n1601) );
  DFFRX1 \CACHE_reg[6][98]  ( .D(n2840), .CK(clk), .RN(n3819), .Q(
        \CACHE[6][98] ), .QN(n1600) );
  DFFRX1 \CACHE_reg[6][97]  ( .D(n2839), .CK(clk), .RN(n3819), .Q(
        \CACHE[6][97] ), .QN(n1599) );
  DFFRX1 \CACHE_reg[6][96]  ( .D(n2838), .CK(clk), .RN(n3819), .Q(
        \CACHE[6][96] ), .QN(n1598) );
  DFFRX1 \CACHE_reg[6][95]  ( .D(n2837), .CK(clk), .RN(n3819), .Q(
        \CACHE[6][95] ), .QN(n1597) );
  DFFRX1 \CACHE_reg[6][94]  ( .D(n2836), .CK(clk), .RN(n3819), .Q(
        \CACHE[6][94] ), .QN(n1596) );
  DFFRX1 \CACHE_reg[6][93]  ( .D(n2835), .CK(clk), .RN(n3819), .Q(
        \CACHE[6][93] ), .QN(n1595) );
  DFFRX1 \CACHE_reg[6][92]  ( .D(n2834), .CK(clk), .RN(n3819), .Q(
        \CACHE[6][92] ), .QN(n1594) );
  DFFRX1 \CACHE_reg[6][91]  ( .D(n2833), .CK(clk), .RN(n3819), .Q(
        \CACHE[6][91] ), .QN(n1593) );
  DFFRX1 \CACHE_reg[6][90]  ( .D(n2832), .CK(clk), .RN(n3819), .Q(
        \CACHE[6][90] ), .QN(n1592) );
  DFFRX1 \CACHE_reg[6][89]  ( .D(n2831), .CK(clk), .RN(n3818), .Q(
        \CACHE[6][89] ), .QN(n1591) );
  DFFRX1 \CACHE_reg[6][88]  ( .D(n2830), .CK(clk), .RN(n3818), .Q(
        \CACHE[6][88] ), .QN(n1590) );
  DFFRX1 \CACHE_reg[6][87]  ( .D(n2829), .CK(clk), .RN(n3818), .Q(
        \CACHE[6][87] ), .QN(n1589) );
  DFFRX1 \CACHE_reg[6][86]  ( .D(n2828), .CK(clk), .RN(n3818), .Q(
        \CACHE[6][86] ), .QN(n1588) );
  DFFRX1 \CACHE_reg[6][85]  ( .D(n2827), .CK(clk), .RN(n3818), .Q(
        \CACHE[6][85] ), .QN(n1587) );
  DFFRX1 \CACHE_reg[6][84]  ( .D(n2826), .CK(clk), .RN(n3818), .Q(
        \CACHE[6][84] ), .QN(n1586) );
  DFFRX1 \CACHE_reg[6][83]  ( .D(n2825), .CK(clk), .RN(n3818), .Q(
        \CACHE[6][83] ), .QN(n1585) );
  DFFRX1 \CACHE_reg[6][82]  ( .D(n2824), .CK(clk), .RN(n3818), .Q(
        \CACHE[6][82] ), .QN(n1584) );
  DFFRX1 \CACHE_reg[6][81]  ( .D(n2823), .CK(clk), .RN(n3818), .Q(
        \CACHE[6][81] ), .QN(n1583) );
  DFFRX1 \CACHE_reg[6][80]  ( .D(n2822), .CK(clk), .RN(n3818), .Q(
        \CACHE[6][80] ), .QN(n1582) );
  DFFRX1 \CACHE_reg[6][79]  ( .D(n2821), .CK(clk), .RN(n3818), .Q(
        \CACHE[6][79] ), .QN(n1581) );
  DFFRX1 \CACHE_reg[6][78]  ( .D(n2820), .CK(clk), .RN(n3818), .Q(
        \CACHE[6][78] ), .QN(n1580) );
  DFFRX1 \CACHE_reg[6][77]  ( .D(n2819), .CK(clk), .RN(n3817), .Q(
        \CACHE[6][77] ), .QN(n1579) );
  DFFRX1 \CACHE_reg[6][76]  ( .D(n2818), .CK(clk), .RN(n3817), .Q(
        \CACHE[6][76] ), .QN(n1578) );
  DFFRX1 \CACHE_reg[6][75]  ( .D(n2817), .CK(clk), .RN(n3817), .Q(
        \CACHE[6][75] ), .QN(n1577) );
  DFFRX1 \CACHE_reg[6][74]  ( .D(n2816), .CK(clk), .RN(n3817), .Q(
        \CACHE[6][74] ), .QN(n1576) );
  DFFRX1 \CACHE_reg[6][73]  ( .D(n2815), .CK(clk), .RN(n3817), .Q(
        \CACHE[6][73] ), .QN(n1575) );
  DFFRX1 \CACHE_reg[6][72]  ( .D(n2814), .CK(clk), .RN(n3817), .Q(
        \CACHE[6][72] ), .QN(n1574) );
  DFFRX1 \CACHE_reg[6][71]  ( .D(n2813), .CK(clk), .RN(n3817), .Q(
        \CACHE[6][71] ), .QN(n1573) );
  DFFRX1 \CACHE_reg[6][70]  ( .D(n2812), .CK(clk), .RN(n3817), .Q(
        \CACHE[6][70] ), .QN(n1572) );
  DFFRX1 \CACHE_reg[6][69]  ( .D(n2811), .CK(clk), .RN(n3817), .Q(
        \CACHE[6][69] ), .QN(n1571) );
  DFFRX1 \CACHE_reg[6][68]  ( .D(n2810), .CK(clk), .RN(n3817), .Q(
        \CACHE[6][68] ), .QN(n1570) );
  DFFRX1 \CACHE_reg[6][67]  ( .D(n2809), .CK(clk), .RN(n3817), .Q(
        \CACHE[6][67] ), .QN(n1569) );
  DFFRX1 \CACHE_reg[6][66]  ( .D(n2808), .CK(clk), .RN(n3817), .Q(
        \CACHE[6][66] ), .QN(n1568) );
  DFFRX1 \CACHE_reg[6][65]  ( .D(n2807), .CK(clk), .RN(n3816), .Q(
        \CACHE[6][65] ), .QN(n1567) );
  DFFRX1 \CACHE_reg[6][64]  ( .D(n2806), .CK(clk), .RN(n3816), .Q(
        \CACHE[6][64] ), .QN(n1566) );
  DFFRX1 \CACHE_reg[6][63]  ( .D(n2805), .CK(clk), .RN(n3816), .Q(
        \CACHE[6][63] ), .QN(n1565) );
  DFFRX1 \CACHE_reg[6][62]  ( .D(n2804), .CK(clk), .RN(n3816), .Q(
        \CACHE[6][62] ), .QN(n1564) );
  DFFRX1 \CACHE_reg[6][61]  ( .D(n2803), .CK(clk), .RN(n3816), .Q(
        \CACHE[6][61] ), .QN(n1563) );
  DFFRX1 \CACHE_reg[6][60]  ( .D(n2802), .CK(clk), .RN(n3816), .Q(
        \CACHE[6][60] ), .QN(n1562) );
  DFFRX1 \CACHE_reg[6][59]  ( .D(n2801), .CK(clk), .RN(n3816), .Q(
        \CACHE[6][59] ), .QN(n1561) );
  DFFRX1 \CACHE_reg[6][58]  ( .D(n2800), .CK(clk), .RN(n3816), .Q(
        \CACHE[6][58] ), .QN(n1560) );
  DFFRX1 \CACHE_reg[6][57]  ( .D(n2799), .CK(clk), .RN(n3816), .Q(
        \CACHE[6][57] ), .QN(n1559) );
  DFFRX1 \CACHE_reg[6][56]  ( .D(n2798), .CK(clk), .RN(n3816), .Q(
        \CACHE[6][56] ), .QN(n1558) );
  DFFRX1 \CACHE_reg[6][55]  ( .D(n2797), .CK(clk), .RN(n3816), .Q(
        \CACHE[6][55] ), .QN(n1557) );
  DFFRX1 \CACHE_reg[6][54]  ( .D(n2796), .CK(clk), .RN(n3816), .Q(
        \CACHE[6][54] ), .QN(n1556) );
  DFFRX1 \CACHE_reg[6][53]  ( .D(n2795), .CK(clk), .RN(n3815), .Q(
        \CACHE[6][53] ), .QN(n1555) );
  DFFRX1 \CACHE_reg[6][52]  ( .D(n2794), .CK(clk), .RN(n3815), .Q(
        \CACHE[6][52] ), .QN(n1554) );
  DFFRX1 \CACHE_reg[6][51]  ( .D(n2793), .CK(clk), .RN(n3815), .Q(
        \CACHE[6][51] ), .QN(n1553) );
  DFFRX1 \CACHE_reg[6][50]  ( .D(n2792), .CK(clk), .RN(n3815), .Q(
        \CACHE[6][50] ), .QN(n1552) );
  DFFRX1 \CACHE_reg[6][49]  ( .D(n2791), .CK(clk), .RN(n3815), .Q(
        \CACHE[6][49] ), .QN(n1551) );
  DFFRX1 \CACHE_reg[6][48]  ( .D(n2790), .CK(clk), .RN(n3815), .Q(
        \CACHE[6][48] ), .QN(n1550) );
  DFFRX1 \CACHE_reg[6][47]  ( .D(n2789), .CK(clk), .RN(n3815), .Q(
        \CACHE[6][47] ), .QN(n1549) );
  DFFRX1 \CACHE_reg[6][46]  ( .D(n2788), .CK(clk), .RN(n3815), .Q(
        \CACHE[6][46] ), .QN(n1548) );
  DFFRX1 \CACHE_reg[6][45]  ( .D(n2787), .CK(clk), .RN(n3815), .Q(
        \CACHE[6][45] ), .QN(n1547) );
  DFFRX1 \CACHE_reg[6][44]  ( .D(n2786), .CK(clk), .RN(n3815), .Q(
        \CACHE[6][44] ), .QN(n1546) );
  DFFRX1 \CACHE_reg[6][43]  ( .D(n2785), .CK(clk), .RN(n3815), .Q(
        \CACHE[6][43] ), .QN(n1545) );
  DFFRX1 \CACHE_reg[6][42]  ( .D(n2784), .CK(clk), .RN(n3815), .Q(
        \CACHE[6][42] ), .QN(n1544) );
  DFFRX1 \CACHE_reg[6][41]  ( .D(n2783), .CK(clk), .RN(n3814), .Q(
        \CACHE[6][41] ), .QN(n1543) );
  DFFRX1 \CACHE_reg[6][40]  ( .D(n2782), .CK(clk), .RN(n3814), .Q(
        \CACHE[6][40] ), .QN(n1542) );
  DFFRX1 \CACHE_reg[6][39]  ( .D(n2781), .CK(clk), .RN(n3814), .Q(
        \CACHE[6][39] ), .QN(n1541) );
  DFFRX1 \CACHE_reg[6][38]  ( .D(n2780), .CK(clk), .RN(n3814), .Q(
        \CACHE[6][38] ), .QN(n1540) );
  DFFRX1 \CACHE_reg[6][37]  ( .D(n2779), .CK(clk), .RN(n3814), .Q(
        \CACHE[6][37] ), .QN(n1539) );
  DFFRX1 \CACHE_reg[6][36]  ( .D(n2778), .CK(clk), .RN(n3814), .Q(
        \CACHE[6][36] ), .QN(n1538) );
  DFFRX1 \CACHE_reg[6][35]  ( .D(n2777), .CK(clk), .RN(n3814), .Q(
        \CACHE[6][35] ), .QN(n1537) );
  DFFRX1 \CACHE_reg[6][34]  ( .D(n2776), .CK(clk), .RN(n3814), .Q(
        \CACHE[6][34] ), .QN(n1536) );
  DFFRX1 \CACHE_reg[6][33]  ( .D(n2775), .CK(clk), .RN(n3814), .Q(
        \CACHE[6][33] ), .QN(n1535) );
  DFFRX1 \CACHE_reg[6][32]  ( .D(n2774), .CK(clk), .RN(n3814), .Q(
        \CACHE[6][32] ), .QN(n1534) );
  DFFRX1 \CACHE_reg[6][31]  ( .D(n2773), .CK(clk), .RN(n3814), .Q(
        \CACHE[6][31] ), .QN(n1533) );
  DFFRX1 \CACHE_reg[6][30]  ( .D(n2772), .CK(clk), .RN(n3814), .Q(
        \CACHE[6][30] ), .QN(n1532) );
  DFFRX1 \CACHE_reg[6][29]  ( .D(n2771), .CK(clk), .RN(n3813), .Q(
        \CACHE[6][29] ), .QN(n1531) );
  DFFRX1 \CACHE_reg[6][28]  ( .D(n2770), .CK(clk), .RN(n3813), .Q(
        \CACHE[6][28] ), .QN(n1530) );
  DFFRX1 \CACHE_reg[6][27]  ( .D(n2769), .CK(clk), .RN(n3813), .Q(
        \CACHE[6][27] ), .QN(n1529) );
  DFFRX1 \CACHE_reg[6][26]  ( .D(n2768), .CK(clk), .RN(n3813), .Q(
        \CACHE[6][26] ), .QN(n1528) );
  DFFRX1 \CACHE_reg[6][25]  ( .D(n2767), .CK(clk), .RN(n3813), .Q(
        \CACHE[6][25] ), .QN(n1527) );
  DFFRX1 \CACHE_reg[6][24]  ( .D(n2766), .CK(clk), .RN(n3813), .Q(
        \CACHE[6][24] ), .QN(n1526) );
  DFFRX1 \CACHE_reg[6][23]  ( .D(n2765), .CK(clk), .RN(n3813), .Q(
        \CACHE[6][23] ), .QN(n1525) );
  DFFRX1 \CACHE_reg[6][22]  ( .D(n2764), .CK(clk), .RN(n3813), .Q(
        \CACHE[6][22] ), .QN(n1524) );
  DFFRX1 \CACHE_reg[6][21]  ( .D(n2763), .CK(clk), .RN(n3813), .Q(
        \CACHE[6][21] ), .QN(n1523) );
  DFFRX1 \CACHE_reg[6][20]  ( .D(n2762), .CK(clk), .RN(n3813), .Q(
        \CACHE[6][20] ), .QN(n1522) );
  DFFRX1 \CACHE_reg[6][19]  ( .D(n2761), .CK(clk), .RN(n3813), .Q(
        \CACHE[6][19] ), .QN(n1521) );
  DFFRX1 \CACHE_reg[6][18]  ( .D(n2760), .CK(clk), .RN(n3813), .Q(
        \CACHE[6][18] ), .QN(n1520) );
  DFFRX1 \CACHE_reg[6][17]  ( .D(n2759), .CK(clk), .RN(n3812), .Q(
        \CACHE[6][17] ), .QN(n1519) );
  DFFRX1 \CACHE_reg[6][16]  ( .D(n2758), .CK(clk), .RN(n3812), .Q(
        \CACHE[6][16] ), .QN(n1518) );
  DFFRX1 \CACHE_reg[6][15]  ( .D(n2757), .CK(clk), .RN(n3812), .Q(
        \CACHE[6][15] ), .QN(n1517) );
  DFFRX1 \CACHE_reg[6][14]  ( .D(n2756), .CK(clk), .RN(n3812), .Q(
        \CACHE[6][14] ), .QN(n1516) );
  DFFRX1 \CACHE_reg[6][13]  ( .D(n2755), .CK(clk), .RN(n3812), .Q(
        \CACHE[6][13] ), .QN(n1515) );
  DFFRX1 \CACHE_reg[6][12]  ( .D(n2754), .CK(clk), .RN(n3812), .Q(
        \CACHE[6][12] ), .QN(n1514) );
  DFFRX1 \CACHE_reg[6][11]  ( .D(n2753), .CK(clk), .RN(n3812), .Q(
        \CACHE[6][11] ), .QN(n1513) );
  DFFRX1 \CACHE_reg[6][10]  ( .D(n2752), .CK(clk), .RN(n3812), .Q(
        \CACHE[6][10] ), .QN(n1512) );
  DFFRX1 \CACHE_reg[6][9]  ( .D(n2751), .CK(clk), .RN(n3812), .Q(\CACHE[6][9] ), .QN(n1511) );
  DFFRX1 \CACHE_reg[6][8]  ( .D(n2750), .CK(clk), .RN(n3812), .Q(\CACHE[6][8] ), .QN(n1510) );
  DFFRX1 \CACHE_reg[6][7]  ( .D(n2749), .CK(clk), .RN(n3812), .Q(\CACHE[6][7] ), .QN(n1509) );
  DFFRX1 \CACHE_reg[6][6]  ( .D(n2748), .CK(clk), .RN(n3812), .Q(\CACHE[6][6] ), .QN(n1508) );
  DFFRX1 \CACHE_reg[6][5]  ( .D(n2747), .CK(clk), .RN(n3811), .Q(\CACHE[6][5] ), .QN(n1507) );
  DFFRX1 \CACHE_reg[6][4]  ( .D(n2746), .CK(clk), .RN(n3811), .Q(\CACHE[6][4] ), .QN(n1506) );
  DFFRX1 \CACHE_reg[6][3]  ( .D(n2745), .CK(clk), .RN(n3811), .Q(\CACHE[6][3] ), .QN(n1505) );
  DFFRX1 \CACHE_reg[6][2]  ( .D(n2744), .CK(clk), .RN(n3811), .Q(\CACHE[6][2] ), .QN(n1504) );
  DFFRX1 \CACHE_reg[6][1]  ( .D(n2743), .CK(clk), .RN(n3811), .Q(\CACHE[6][1] ), .QN(n1503) );
  DFFRX1 \CACHE_reg[6][0]  ( .D(n2742), .CK(clk), .RN(n3811), .Q(\CACHE[6][0] ), .QN(n1502) );
  DFFRX1 \CACHE_reg[2][118]  ( .D(n2240), .CK(clk), .RN(n3769), .Q(
        \CACHE[2][118] ), .QN(n1000) );
  DFFRX1 \CACHE_reg[2][117]  ( .D(n2239), .CK(clk), .RN(n3769), .Q(
        \CACHE[2][117] ), .QN(n999) );
  DFFRX1 \CACHE_reg[2][116]  ( .D(n2238), .CK(clk), .RN(n3769), .Q(
        \CACHE[2][116] ), .QN(n998) );
  DFFRX1 \CACHE_reg[2][115]  ( .D(n2237), .CK(clk), .RN(n3769), .Q(
        \CACHE[2][115] ), .QN(n997) );
  DFFRX1 \CACHE_reg[2][114]  ( .D(n2236), .CK(clk), .RN(n3769), .Q(
        \CACHE[2][114] ), .QN(n996) );
  DFFRX1 \CACHE_reg[2][113]  ( .D(n2235), .CK(clk), .RN(n3769), .Q(
        \CACHE[2][113] ), .QN(n995) );
  DFFRX1 \CACHE_reg[2][112]  ( .D(n2234), .CK(clk), .RN(n3769), .Q(
        \CACHE[2][112] ), .QN(n994) );
  DFFRX1 \CACHE_reg[2][111]  ( .D(n2233), .CK(clk), .RN(n3769), .Q(
        \CACHE[2][111] ), .QN(n993) );
  DFFRX1 \CACHE_reg[2][110]  ( .D(n2232), .CK(clk), .RN(n3769), .Q(
        \CACHE[2][110] ), .QN(n992) );
  DFFRX1 \CACHE_reg[2][109]  ( .D(n2231), .CK(clk), .RN(n3768), .Q(
        \CACHE[2][109] ), .QN(n991) );
  DFFRX1 \CACHE_reg[2][108]  ( .D(n2230), .CK(clk), .RN(n3768), .Q(
        \CACHE[2][108] ), .QN(n990) );
  DFFRX1 \CACHE_reg[2][107]  ( .D(n2229), .CK(clk), .RN(n3768), .Q(
        \CACHE[2][107] ), .QN(n989) );
  DFFRX1 \CACHE_reg[2][106]  ( .D(n2228), .CK(clk), .RN(n3768), .Q(
        \CACHE[2][106] ), .QN(n988) );
  DFFRX1 \CACHE_reg[2][105]  ( .D(n2227), .CK(clk), .RN(n3768), .Q(
        \CACHE[2][105] ), .QN(n987) );
  DFFRX1 \CACHE_reg[2][104]  ( .D(n2226), .CK(clk), .RN(n3768), .Q(
        \CACHE[2][104] ), .QN(n986) );
  DFFRX1 \CACHE_reg[2][103]  ( .D(n2225), .CK(clk), .RN(n3768), .Q(
        \CACHE[2][103] ), .QN(n985) );
  DFFRX1 \CACHE_reg[2][102]  ( .D(n2224), .CK(clk), .RN(n3768), .Q(
        \CACHE[2][102] ), .QN(n984) );
  DFFRX1 \CACHE_reg[2][101]  ( .D(n2223), .CK(clk), .RN(n3768), .Q(
        \CACHE[2][101] ), .QN(n983) );
  DFFRX1 \CACHE_reg[2][100]  ( .D(n2222), .CK(clk), .RN(n3768), .Q(
        \CACHE[2][100] ), .QN(n982) );
  DFFRX1 \CACHE_reg[2][99]  ( .D(n2221), .CK(clk), .RN(n3768), .Q(
        \CACHE[2][99] ), .QN(n981) );
  DFFRX1 \CACHE_reg[2][98]  ( .D(n2220), .CK(clk), .RN(n3768), .Q(
        \CACHE[2][98] ), .QN(n980) );
  DFFRX1 \CACHE_reg[2][97]  ( .D(n2219), .CK(clk), .RN(n3767), .Q(
        \CACHE[2][97] ), .QN(n979) );
  DFFRX1 \CACHE_reg[2][96]  ( .D(n2218), .CK(clk), .RN(n3767), .Q(
        \CACHE[2][96] ), .QN(n978) );
  DFFRX1 \CACHE_reg[2][95]  ( .D(n2217), .CK(clk), .RN(n3767), .Q(
        \CACHE[2][95] ), .QN(n977) );
  DFFRX1 \CACHE_reg[2][94]  ( .D(n2216), .CK(clk), .RN(n3767), .Q(
        \CACHE[2][94] ), .QN(n976) );
  DFFRX1 \CACHE_reg[2][93]  ( .D(n2215), .CK(clk), .RN(n3767), .Q(
        \CACHE[2][93] ), .QN(n975) );
  DFFRX1 \CACHE_reg[2][92]  ( .D(n2214), .CK(clk), .RN(n3767), .Q(
        \CACHE[2][92] ), .QN(n974) );
  DFFRX1 \CACHE_reg[2][91]  ( .D(n2213), .CK(clk), .RN(n3767), .Q(
        \CACHE[2][91] ), .QN(n973) );
  DFFRX1 \CACHE_reg[2][90]  ( .D(n2212), .CK(clk), .RN(n3767), .Q(
        \CACHE[2][90] ), .QN(n972) );
  DFFRX1 \CACHE_reg[2][89]  ( .D(n2211), .CK(clk), .RN(n3767), .Q(
        \CACHE[2][89] ), .QN(n971) );
  DFFRX1 \CACHE_reg[2][88]  ( .D(n2210), .CK(clk), .RN(n3767), .Q(
        \CACHE[2][88] ), .QN(n970) );
  DFFRX1 \CACHE_reg[2][87]  ( .D(n2209), .CK(clk), .RN(n3767), .Q(
        \CACHE[2][87] ), .QN(n969) );
  DFFRX1 \CACHE_reg[2][86]  ( .D(n2208), .CK(clk), .RN(n3767), .Q(
        \CACHE[2][86] ), .QN(n968) );
  DFFRX1 \CACHE_reg[2][85]  ( .D(n2207), .CK(clk), .RN(n3766), .Q(
        \CACHE[2][85] ), .QN(n967) );
  DFFRX1 \CACHE_reg[2][84]  ( .D(n2206), .CK(clk), .RN(n3766), .Q(
        \CACHE[2][84] ), .QN(n966) );
  DFFRX1 \CACHE_reg[2][83]  ( .D(n2205), .CK(clk), .RN(n3766), .Q(
        \CACHE[2][83] ), .QN(n965) );
  DFFRX1 \CACHE_reg[2][82]  ( .D(n2204), .CK(clk), .RN(n3766), .Q(
        \CACHE[2][82] ), .QN(n964) );
  DFFRX1 \CACHE_reg[2][81]  ( .D(n2203), .CK(clk), .RN(n3766), .Q(
        \CACHE[2][81] ), .QN(n963) );
  DFFRX1 \CACHE_reg[2][80]  ( .D(n2202), .CK(clk), .RN(n3766), .Q(
        \CACHE[2][80] ), .QN(n962) );
  DFFRX1 \CACHE_reg[2][79]  ( .D(n2201), .CK(clk), .RN(n3766), .Q(
        \CACHE[2][79] ), .QN(n961) );
  DFFRX1 \CACHE_reg[2][78]  ( .D(n2200), .CK(clk), .RN(n3766), .Q(
        \CACHE[2][78] ), .QN(n960) );
  DFFRX1 \CACHE_reg[2][77]  ( .D(n2199), .CK(clk), .RN(n3766), .Q(
        \CACHE[2][77] ), .QN(n959) );
  DFFRX1 \CACHE_reg[2][76]  ( .D(n2198), .CK(clk), .RN(n3766), .Q(
        \CACHE[2][76] ), .QN(n958) );
  DFFRX1 \CACHE_reg[2][75]  ( .D(n2197), .CK(clk), .RN(n3766), .Q(
        \CACHE[2][75] ), .QN(n957) );
  DFFRX1 \CACHE_reg[2][74]  ( .D(n2196), .CK(clk), .RN(n3766), .Q(
        \CACHE[2][74] ), .QN(n956) );
  DFFRX1 \CACHE_reg[2][73]  ( .D(n2195), .CK(clk), .RN(n3765), .Q(
        \CACHE[2][73] ), .QN(n955) );
  DFFRX1 \CACHE_reg[2][72]  ( .D(n2194), .CK(clk), .RN(n3765), .Q(
        \CACHE[2][72] ), .QN(n954) );
  DFFRX1 \CACHE_reg[2][71]  ( .D(n2193), .CK(clk), .RN(n3765), .Q(
        \CACHE[2][71] ), .QN(n953) );
  DFFRX1 \CACHE_reg[2][70]  ( .D(n2192), .CK(clk), .RN(n3765), .Q(
        \CACHE[2][70] ), .QN(n952) );
  DFFRX1 \CACHE_reg[2][69]  ( .D(n2191), .CK(clk), .RN(n3765), .Q(
        \CACHE[2][69] ), .QN(n951) );
  DFFRX1 \CACHE_reg[2][68]  ( .D(n2190), .CK(clk), .RN(n3765), .Q(
        \CACHE[2][68] ), .QN(n950) );
  DFFRX1 \CACHE_reg[2][67]  ( .D(n2189), .CK(clk), .RN(n3765), .Q(
        \CACHE[2][67] ), .QN(n949) );
  DFFRX1 \CACHE_reg[2][66]  ( .D(n2188), .CK(clk), .RN(n3765), .Q(
        \CACHE[2][66] ), .QN(n948) );
  DFFRX1 \CACHE_reg[2][65]  ( .D(n2187), .CK(clk), .RN(n3765), .Q(
        \CACHE[2][65] ), .QN(n947) );
  DFFRX1 \CACHE_reg[2][64]  ( .D(n2186), .CK(clk), .RN(n3765), .Q(
        \CACHE[2][64] ), .QN(n946) );
  DFFRX1 \CACHE_reg[2][63]  ( .D(n2185), .CK(clk), .RN(n3765), .Q(
        \CACHE[2][63] ), .QN(n945) );
  DFFRX1 \CACHE_reg[2][62]  ( .D(n2184), .CK(clk), .RN(n3765), .Q(
        \CACHE[2][62] ), .QN(n944) );
  DFFRX1 \CACHE_reg[2][61]  ( .D(n2183), .CK(clk), .RN(n3764), .Q(
        \CACHE[2][61] ), .QN(n943) );
  DFFRX1 \CACHE_reg[2][60]  ( .D(n2182), .CK(clk), .RN(n3764), .Q(
        \CACHE[2][60] ), .QN(n942) );
  DFFRX1 \CACHE_reg[2][59]  ( .D(n2181), .CK(clk), .RN(n3764), .Q(
        \CACHE[2][59] ), .QN(n941) );
  DFFRX1 \CACHE_reg[2][58]  ( .D(n2180), .CK(clk), .RN(n3764), .Q(
        \CACHE[2][58] ), .QN(n940) );
  DFFRX1 \CACHE_reg[2][57]  ( .D(n2179), .CK(clk), .RN(n3764), .Q(
        \CACHE[2][57] ), .QN(n939) );
  DFFRX1 \CACHE_reg[2][56]  ( .D(n2178), .CK(clk), .RN(n3764), .Q(
        \CACHE[2][56] ), .QN(n938) );
  DFFRX1 \CACHE_reg[2][55]  ( .D(n2177), .CK(clk), .RN(n3764), .Q(
        \CACHE[2][55] ), .QN(n937) );
  DFFRX1 \CACHE_reg[2][54]  ( .D(n2176), .CK(clk), .RN(n3764), .Q(
        \CACHE[2][54] ), .QN(n936) );
  DFFRX1 \CACHE_reg[2][53]  ( .D(n2175), .CK(clk), .RN(n3764), .Q(
        \CACHE[2][53] ), .QN(n935) );
  DFFRX1 \CACHE_reg[2][52]  ( .D(n2174), .CK(clk), .RN(n3764), .Q(
        \CACHE[2][52] ), .QN(n934) );
  DFFRX1 \CACHE_reg[2][51]  ( .D(n2173), .CK(clk), .RN(n3764), .Q(
        \CACHE[2][51] ), .QN(n933) );
  DFFRX1 \CACHE_reg[2][50]  ( .D(n2172), .CK(clk), .RN(n3764), .Q(
        \CACHE[2][50] ), .QN(n932) );
  DFFRX1 \CACHE_reg[2][49]  ( .D(n2171), .CK(clk), .RN(n3763), .Q(
        \CACHE[2][49] ), .QN(n931) );
  DFFRX1 \CACHE_reg[2][48]  ( .D(n2170), .CK(clk), .RN(n3763), .Q(
        \CACHE[2][48] ), .QN(n930) );
  DFFRX1 \CACHE_reg[2][47]  ( .D(n2169), .CK(clk), .RN(n3763), .Q(
        \CACHE[2][47] ), .QN(n929) );
  DFFRX1 \CACHE_reg[2][46]  ( .D(n2168), .CK(clk), .RN(n3763), .Q(
        \CACHE[2][46] ), .QN(n928) );
  DFFRX1 \CACHE_reg[2][45]  ( .D(n2167), .CK(clk), .RN(n3763), .Q(
        \CACHE[2][45] ), .QN(n927) );
  DFFRX1 \CACHE_reg[2][44]  ( .D(n2166), .CK(clk), .RN(n3763), .Q(
        \CACHE[2][44] ), .QN(n926) );
  DFFRX1 \CACHE_reg[2][43]  ( .D(n2165), .CK(clk), .RN(n3763), .Q(
        \CACHE[2][43] ), .QN(n925) );
  DFFRX1 \CACHE_reg[2][42]  ( .D(n2164), .CK(clk), .RN(n3763), .Q(
        \CACHE[2][42] ), .QN(n924) );
  DFFRX1 \CACHE_reg[2][41]  ( .D(n2163), .CK(clk), .RN(n3763), .Q(
        \CACHE[2][41] ), .QN(n923) );
  DFFRX1 \CACHE_reg[2][40]  ( .D(n2162), .CK(clk), .RN(n3763), .Q(
        \CACHE[2][40] ), .QN(n922) );
  DFFRX1 \CACHE_reg[2][39]  ( .D(n2161), .CK(clk), .RN(n3763), .Q(
        \CACHE[2][39] ), .QN(n921) );
  DFFRX1 \CACHE_reg[2][38]  ( .D(n2160), .CK(clk), .RN(n3763), .Q(
        \CACHE[2][38] ), .QN(n920) );
  DFFRX1 \CACHE_reg[2][37]  ( .D(n2159), .CK(clk), .RN(n3762), .Q(
        \CACHE[2][37] ), .QN(n919) );
  DFFRX1 \CACHE_reg[2][36]  ( .D(n2158), .CK(clk), .RN(n3762), .Q(
        \CACHE[2][36] ), .QN(n918) );
  DFFRX1 \CACHE_reg[2][35]  ( .D(n2157), .CK(clk), .RN(n3762), .Q(
        \CACHE[2][35] ), .QN(n917) );
  DFFRX1 \CACHE_reg[2][34]  ( .D(n2156), .CK(clk), .RN(n3762), .Q(
        \CACHE[2][34] ), .QN(n916) );
  DFFRX1 \CACHE_reg[2][33]  ( .D(n2155), .CK(clk), .RN(n3762), .Q(
        \CACHE[2][33] ), .QN(n915) );
  DFFRX1 \CACHE_reg[2][32]  ( .D(n2154), .CK(clk), .RN(n3762), .Q(
        \CACHE[2][32] ), .QN(n914) );
  DFFRX1 \CACHE_reg[2][31]  ( .D(n2153), .CK(clk), .RN(n3762), .Q(
        \CACHE[2][31] ), .QN(n913) );
  DFFRX1 \CACHE_reg[2][30]  ( .D(n2152), .CK(clk), .RN(n3762), .Q(
        \CACHE[2][30] ), .QN(n912) );
  DFFRX1 \CACHE_reg[2][29]  ( .D(n2151), .CK(clk), .RN(n3762), .Q(
        \CACHE[2][29] ), .QN(n911) );
  DFFRX1 \CACHE_reg[2][28]  ( .D(n2150), .CK(clk), .RN(n3762), .Q(
        \CACHE[2][28] ), .QN(n910) );
  DFFRX1 \CACHE_reg[2][27]  ( .D(n2149), .CK(clk), .RN(n3762), .Q(
        \CACHE[2][27] ), .QN(n909) );
  DFFRX1 \CACHE_reg[2][26]  ( .D(n2148), .CK(clk), .RN(n3762), .Q(
        \CACHE[2][26] ), .QN(n908) );
  DFFRX1 \CACHE_reg[2][25]  ( .D(n2147), .CK(clk), .RN(n3761), .Q(
        \CACHE[2][25] ), .QN(n907) );
  DFFRX1 \CACHE_reg[2][24]  ( .D(n2146), .CK(clk), .RN(n3761), .Q(
        \CACHE[2][24] ), .QN(n906) );
  DFFRX1 \CACHE_reg[2][23]  ( .D(n2145), .CK(clk), .RN(n3761), .Q(
        \CACHE[2][23] ), .QN(n905) );
  DFFRX1 \CACHE_reg[2][22]  ( .D(n2144), .CK(clk), .RN(n3761), .Q(
        \CACHE[2][22] ), .QN(n904) );
  DFFRX1 \CACHE_reg[2][21]  ( .D(n2143), .CK(clk), .RN(n3761), .Q(
        \CACHE[2][21] ), .QN(n903) );
  DFFRX1 \CACHE_reg[2][20]  ( .D(n2142), .CK(clk), .RN(n3761), .Q(
        \CACHE[2][20] ), .QN(n902) );
  DFFRX1 \CACHE_reg[2][19]  ( .D(n2141), .CK(clk), .RN(n3761), .Q(
        \CACHE[2][19] ), .QN(n901) );
  DFFRX1 \CACHE_reg[2][18]  ( .D(n2140), .CK(clk), .RN(n3761), .Q(
        \CACHE[2][18] ), .QN(n900) );
  DFFRX1 \CACHE_reg[2][17]  ( .D(n2139), .CK(clk), .RN(n3761), .Q(
        \CACHE[2][17] ), .QN(n899) );
  DFFRX1 \CACHE_reg[2][16]  ( .D(n2138), .CK(clk), .RN(n3761), .Q(
        \CACHE[2][16] ), .QN(n898) );
  DFFRX1 \CACHE_reg[2][15]  ( .D(n2137), .CK(clk), .RN(n3761), .Q(
        \CACHE[2][15] ), .QN(n897) );
  DFFRX1 \CACHE_reg[2][14]  ( .D(n2136), .CK(clk), .RN(n3761), .Q(
        \CACHE[2][14] ), .QN(n896) );
  DFFRX1 \CACHE_reg[2][13]  ( .D(n2135), .CK(clk), .RN(n3760), .Q(
        \CACHE[2][13] ), .QN(n895) );
  DFFRX1 \CACHE_reg[2][12]  ( .D(n2134), .CK(clk), .RN(n3760), .Q(
        \CACHE[2][12] ), .QN(n894) );
  DFFRX1 \CACHE_reg[2][11]  ( .D(n2133), .CK(clk), .RN(n3760), .Q(
        \CACHE[2][11] ), .QN(n893) );
  DFFRX1 \CACHE_reg[2][10]  ( .D(n2132), .CK(clk), .RN(n3760), .Q(
        \CACHE[2][10] ), .QN(n892) );
  DFFRX1 \CACHE_reg[2][9]  ( .D(n2131), .CK(clk), .RN(n3760), .Q(\CACHE[2][9] ), .QN(n891) );
  DFFRX1 \CACHE_reg[2][8]  ( .D(n2130), .CK(clk), .RN(n3760), .Q(\CACHE[2][8] ), .QN(n890) );
  DFFRX1 \CACHE_reg[2][7]  ( .D(n2129), .CK(clk), .RN(n3760), .Q(\CACHE[2][7] ), .QN(n889) );
  DFFRX1 \CACHE_reg[2][6]  ( .D(n2128), .CK(clk), .RN(n3760), .Q(\CACHE[2][6] ), .QN(n888) );
  DFFRX1 \CACHE_reg[2][5]  ( .D(n2127), .CK(clk), .RN(n3760), .Q(\CACHE[2][5] ), .QN(n887) );
  DFFRX1 \CACHE_reg[2][4]  ( .D(n2126), .CK(clk), .RN(n3760), .Q(\CACHE[2][4] ), .QN(n886) );
  DFFRX1 \CACHE_reg[2][3]  ( .D(n2125), .CK(clk), .RN(n3760), .Q(\CACHE[2][3] ), .QN(n885) );
  DFFRX1 \CACHE_reg[2][2]  ( .D(n2124), .CK(clk), .RN(n3760), .Q(\CACHE[2][2] ), .QN(n884) );
  DFFRX1 \CACHE_reg[2][0]  ( .D(n2122), .CK(clk), .RN(n3759), .Q(\CACHE[2][0] ), .QN(n882) );
  DFFRX1 \CACHE_reg[7][154]  ( .D(n3052), .CK(clk), .RN(n3837), .QN(n1811) );
  DFFRX1 \CACHE_reg[7][153]  ( .D(n3050), .CK(clk), .RN(n3837), .Q(
        \CACHE[7][153] ), .QN(n1810) );
  DFFRX1 \CACHE_reg[7][152]  ( .D(n3049), .CK(clk), .RN(n3837), .QN(n1809) );
  DFFRX1 \CACHE_reg[7][151]  ( .D(n3048), .CK(clk), .RN(n3837), .QN(n1808) );
  DFFRX1 \CACHE_reg[7][150]  ( .D(n3047), .CK(clk), .RN(n3836), .QN(n1807) );
  DFFRX1 \CACHE_reg[7][149]  ( .D(n3046), .CK(clk), .RN(n3836), .Q(
        \CACHE[7][149] ), .QN(n1806) );
  DFFRX1 \CACHE_reg[7][148]  ( .D(n3045), .CK(clk), .RN(n3836), .Q(
        \CACHE[7][148] ), .QN(n1805) );
  DFFRX1 \CACHE_reg[7][147]  ( .D(n3044), .CK(clk), .RN(n3836), .QN(n1804) );
  DFFRX1 \CACHE_reg[7][146]  ( .D(n3043), .CK(clk), .RN(n3836), .QN(n1803) );
  DFFRX1 \CACHE_reg[7][145]  ( .D(n3042), .CK(clk), .RN(n3836), .QN(n1802) );
  DFFRX1 \CACHE_reg[7][144]  ( .D(n3041), .CK(clk), .RN(n3836), .QN(n1801) );
  DFFRX1 \CACHE_reg[7][143]  ( .D(n3040), .CK(clk), .RN(n3836), .Q(
        \CACHE[7][143] ), .QN(n1800) );
  DFFRX1 \CACHE_reg[7][142]  ( .D(n3039), .CK(clk), .RN(n3836), .Q(
        \CACHE[7][142] ), .QN(n1799) );
  DFFRX1 \CACHE_reg[7][141]  ( .D(n3038), .CK(clk), .RN(n3836), .Q(
        \CACHE[7][141] ), .QN(n1798) );
  DFFRX1 \CACHE_reg[7][140]  ( .D(n3037), .CK(clk), .RN(n3836), .QN(n1797) );
  DFFRX1 \CACHE_reg[7][139]  ( .D(n3036), .CK(clk), .RN(n3836), .Q(
        \CACHE[7][139] ), .QN(n1796) );
  DFFRX1 \CACHE_reg[7][138]  ( .D(n3035), .CK(clk), .RN(n3835), .Q(
        \CACHE[7][138] ), .QN(n1795) );
  DFFRX1 \CACHE_reg[7][137]  ( .D(n3034), .CK(clk), .RN(n3835), .Q(
        \CACHE[7][137] ), .QN(n1794) );
  DFFRX1 \CACHE_reg[7][136]  ( .D(n3033), .CK(clk), .RN(n3835), .Q(
        \CACHE[7][136] ), .QN(n1793) );
  DFFRX1 \CACHE_reg[7][135]  ( .D(n3032), .CK(clk), .RN(n3835), .QN(n1792) );
  DFFRX1 \CACHE_reg[7][134]  ( .D(n3031), .CK(clk), .RN(n3835), .QN(n1791) );
  DFFRX1 \CACHE_reg[7][133]  ( .D(n3030), .CK(clk), .RN(n3835), .QN(n1790) );
  DFFRX1 \CACHE_reg[7][132]  ( .D(n3029), .CK(clk), .RN(n3835), .Q(
        \CACHE[7][132] ), .QN(n1789) );
  DFFRX1 \CACHE_reg[7][131]  ( .D(n3028), .CK(clk), .RN(n3835), .Q(
        \CACHE[7][131] ), .QN(n1788) );
  DFFRX1 \CACHE_reg[7][130]  ( .D(n3027), .CK(clk), .RN(n3835), .QN(n1787) );
  DFFRX1 \CACHE_reg[7][129]  ( .D(n3026), .CK(clk), .RN(n3835), .Q(
        \CACHE[7][129] ), .QN(n1786) );
  DFFRX1 \CACHE_reg[7][128]  ( .D(n3025), .CK(clk), .RN(n3835), .Q(
        \CACHE[7][128] ), .QN(n1785) );
  DFFRX1 \CACHE_reg[3][154]  ( .D(n2431), .CK(clk), .RN(n3785), .QN(n1191) );
  DFFRX1 \CACHE_reg[3][153]  ( .D(n2430), .CK(clk), .RN(n3785), .Q(
        \CACHE[3][153] ), .QN(n1190) );
  DFFRX1 \CACHE_reg[3][152]  ( .D(n2429), .CK(clk), .RN(n3785), .QN(n1189) );
  DFFRX1 \CACHE_reg[3][151]  ( .D(n2428), .CK(clk), .RN(n3785), .QN(n1188) );
  DFFRX1 \CACHE_reg[3][150]  ( .D(n2427), .CK(clk), .RN(n3785), .QN(n1187) );
  DFFRX1 \CACHE_reg[3][149]  ( .D(n2426), .CK(clk), .RN(n3785), .Q(
        \CACHE[3][149] ), .QN(n1186) );
  DFFRX1 \CACHE_reg[3][148]  ( .D(n2425), .CK(clk), .RN(n3785), .Q(
        \CACHE[3][148] ), .QN(n1185) );
  DFFRX1 \CACHE_reg[3][147]  ( .D(n2424), .CK(clk), .RN(n3785), .QN(n1184) );
  DFFRX1 \CACHE_reg[3][146]  ( .D(n2423), .CK(clk), .RN(n3784), .QN(n1183) );
  DFFRX1 \CACHE_reg[3][145]  ( .D(n2422), .CK(clk), .RN(n3784), .QN(n1182) );
  DFFRX1 \CACHE_reg[3][144]  ( .D(n2421), .CK(clk), .RN(n3784), .QN(n1181) );
  DFFRX1 \CACHE_reg[3][143]  ( .D(n2420), .CK(clk), .RN(n3784), .Q(
        \CACHE[3][143] ), .QN(n1180) );
  DFFRX1 \CACHE_reg[3][142]  ( .D(n2419), .CK(clk), .RN(n3784), .Q(
        \CACHE[3][142] ), .QN(n1179) );
  DFFRX1 \CACHE_reg[3][141]  ( .D(n2418), .CK(clk), .RN(n3784), .Q(
        \CACHE[3][141] ), .QN(n1178) );
  DFFRX1 \CACHE_reg[3][140]  ( .D(n2417), .CK(clk), .RN(n3784), .QN(n1177) );
  DFFRX1 \CACHE_reg[3][139]  ( .D(n2416), .CK(clk), .RN(n3784), .Q(
        \CACHE[3][139] ), .QN(n1176) );
  DFFRX1 \CACHE_reg[3][138]  ( .D(n2415), .CK(clk), .RN(n3784), .Q(
        \CACHE[3][138] ), .QN(n1175) );
  DFFRX1 \CACHE_reg[3][137]  ( .D(n2414), .CK(clk), .RN(n3784), .Q(
        \CACHE[3][137] ), .QN(n1174) );
  DFFRX1 \CACHE_reg[3][136]  ( .D(n2413), .CK(clk), .RN(n3784), .Q(
        \CACHE[3][136] ), .QN(n1173) );
  DFFRX1 \CACHE_reg[3][135]  ( .D(n2412), .CK(clk), .RN(n3784), .Q(
        \CACHE[3][135] ), .QN(n1172) );
  DFFRX1 \CACHE_reg[3][134]  ( .D(n2411), .CK(clk), .RN(n3783), .QN(n1171) );
  DFFRX1 \CACHE_reg[3][133]  ( .D(n2410), .CK(clk), .RN(n3783), .QN(n1170) );
  DFFRX1 \CACHE_reg[3][132]  ( .D(n2409), .CK(clk), .RN(n3783), .Q(
        \CACHE[3][132] ), .QN(n1169) );
  DFFRX1 \CACHE_reg[3][131]  ( .D(n2408), .CK(clk), .RN(n3783), .Q(
        \CACHE[3][131] ), .QN(n1168) );
  DFFRX1 \CACHE_reg[3][130]  ( .D(n2407), .CK(clk), .RN(n3783), .QN(n1167) );
  DFFRX1 \CACHE_reg[3][129]  ( .D(n2406), .CK(clk), .RN(n3783), .Q(
        \CACHE[3][129] ), .QN(n1166) );
  DFFRX1 \CACHE_reg[3][128]  ( .D(n2405), .CK(clk), .RN(n3783), .Q(
        \CACHE[3][128] ), .QN(n1165) );
  DFFRX1 \CACHE_reg[5][154]  ( .D(n2741), .CK(clk), .RN(n3811), .QN(n1501) );
  DFFRX1 \CACHE_reg[5][153]  ( .D(n2740), .CK(clk), .RN(n3811), .Q(
        \CACHE[5][153] ), .QN(n1500) );
  DFFRX1 \CACHE_reg[5][152]  ( .D(n2739), .CK(clk), .RN(n3811), .QN(n1499) );
  DFFRX1 \CACHE_reg[5][151]  ( .D(n2738), .CK(clk), .RN(n3811), .QN(n1498) );
  DFFRX1 \CACHE_reg[5][150]  ( .D(n2737), .CK(clk), .RN(n3811), .QN(n1497) );
  DFFRX1 \CACHE_reg[5][149]  ( .D(n2736), .CK(clk), .RN(n3811), .Q(
        \CACHE[5][149] ), .QN(n1496) );
  DFFRX1 \CACHE_reg[5][148]  ( .D(n2735), .CK(clk), .RN(n3810), .Q(
        \CACHE[5][148] ), .QN(n1495) );
  DFFRX1 \CACHE_reg[5][147]  ( .D(n2734), .CK(clk), .RN(n3810), .QN(n1494) );
  DFFRX1 \CACHE_reg[5][146]  ( .D(n2733), .CK(clk), .RN(n3810), .QN(n1493) );
  DFFRX1 \CACHE_reg[5][145]  ( .D(n2732), .CK(clk), .RN(n3810), .QN(n1492) );
  DFFRX1 \CACHE_reg[5][144]  ( .D(n2731), .CK(clk), .RN(n3810), .QN(n1491) );
  DFFRX1 \CACHE_reg[5][143]  ( .D(n2730), .CK(clk), .RN(n3810), .Q(
        \CACHE[5][143] ), .QN(n1490) );
  DFFRX1 \CACHE_reg[5][142]  ( .D(n2729), .CK(clk), .RN(n3810), .Q(
        \CACHE[5][142] ), .QN(n1489) );
  DFFRX1 \CACHE_reg[5][141]  ( .D(n2728), .CK(clk), .RN(n3810), .Q(
        \CACHE[5][141] ), .QN(n1488) );
  DFFRX1 \CACHE_reg[5][140]  ( .D(n2727), .CK(clk), .RN(n3810), .QN(n1487) );
  DFFRX1 \CACHE_reg[5][139]  ( .D(n2726), .CK(clk), .RN(n3810), .Q(
        \CACHE[5][139] ), .QN(n1486) );
  DFFRX1 \CACHE_reg[5][138]  ( .D(n2725), .CK(clk), .RN(n3810), .Q(
        \CACHE[5][138] ), .QN(n1485) );
  DFFRX1 \CACHE_reg[5][137]  ( .D(n2724), .CK(clk), .RN(n3810), .Q(
        \CACHE[5][137] ), .QN(n1484) );
  DFFRX1 \CACHE_reg[5][136]  ( .D(n2723), .CK(clk), .RN(n3809), .Q(
        \CACHE[5][136] ), .QN(n1483) );
  DFFRX1 \CACHE_reg[5][135]  ( .D(n2722), .CK(clk), .RN(n3809), .QN(n1482) );
  DFFRX1 \CACHE_reg[5][134]  ( .D(n2721), .CK(clk), .RN(n3809), .QN(n1481) );
  DFFRX1 \CACHE_reg[5][133]  ( .D(n2720), .CK(clk), .RN(n3809), .QN(n1480) );
  DFFRX1 \CACHE_reg[5][132]  ( .D(n2719), .CK(clk), .RN(n3809), .Q(
        \CACHE[5][132] ), .QN(n1479) );
  DFFRX1 \CACHE_reg[5][131]  ( .D(n2718), .CK(clk), .RN(n3809), .Q(
        \CACHE[5][131] ), .QN(n1478) );
  DFFRX1 \CACHE_reg[5][130]  ( .D(n2717), .CK(clk), .RN(n3809), .QN(n1477) );
  DFFRX1 \CACHE_reg[5][129]  ( .D(n2716), .CK(clk), .RN(n3809), .Q(
        \CACHE[5][129] ), .QN(n1476) );
  DFFRX1 \CACHE_reg[5][128]  ( .D(n2715), .CK(clk), .RN(n3809), .Q(
        \CACHE[5][128] ), .QN(n1475) );
  DFFRX1 \CACHE_reg[1][154]  ( .D(n2121), .CK(clk), .RN(n3759), .QN(n881) );
  DFFRX1 \CACHE_reg[1][153]  ( .D(n2120), .CK(clk), .RN(n3759), .Q(
        \CACHE[1][153] ), .QN(n880) );
  DFFRX1 \CACHE_reg[1][152]  ( .D(n2119), .CK(clk), .RN(n3759), .QN(n879) );
  DFFRX1 \CACHE_reg[1][151]  ( .D(n2118), .CK(clk), .RN(n3759), .QN(n878) );
  DFFRX1 \CACHE_reg[1][150]  ( .D(n2117), .CK(clk), .RN(n3759), .QN(n877) );
  DFFRX1 \CACHE_reg[1][149]  ( .D(n2116), .CK(clk), .RN(n3759), .Q(
        \CACHE[1][149] ), .QN(n876) );
  DFFRX1 \CACHE_reg[1][148]  ( .D(n2115), .CK(clk), .RN(n3759), .Q(
        \CACHE[1][148] ), .QN(n875) );
  DFFRX1 \CACHE_reg[1][147]  ( .D(n2114), .CK(clk), .RN(n3759), .QN(n874) );
  DFFRX1 \CACHE_reg[1][146]  ( .D(n2113), .CK(clk), .RN(n3759), .QN(n873) );
  DFFRX1 \CACHE_reg[1][145]  ( .D(n2112), .CK(clk), .RN(n3759), .QN(n872) );
  DFFRX1 \CACHE_reg[1][144]  ( .D(n2111), .CK(clk), .RN(n3758), .QN(n871) );
  DFFRX1 \CACHE_reg[1][143]  ( .D(n2110), .CK(clk), .RN(n3758), .Q(
        \CACHE[1][143] ), .QN(n870) );
  DFFRX1 \CACHE_reg[1][142]  ( .D(n2109), .CK(clk), .RN(n3758), .Q(
        \CACHE[1][142] ), .QN(n869) );
  DFFRX1 \CACHE_reg[1][141]  ( .D(n2108), .CK(clk), .RN(n3758), .Q(
        \CACHE[1][141] ), .QN(n868) );
  DFFRX1 \CACHE_reg[1][140]  ( .D(n2107), .CK(clk), .RN(n3758), .QN(n867) );
  DFFRX1 \CACHE_reg[1][139]  ( .D(n2106), .CK(clk), .RN(n3758), .Q(
        \CACHE[1][139] ), .QN(n866) );
  DFFRX1 \CACHE_reg[1][138]  ( .D(n2105), .CK(clk), .RN(n3758), .Q(
        \CACHE[1][138] ), .QN(n865) );
  DFFRX1 \CACHE_reg[1][137]  ( .D(n2104), .CK(clk), .RN(n3758), .Q(
        \CACHE[1][137] ), .QN(n864) );
  DFFRX1 \CACHE_reg[1][136]  ( .D(n2103), .CK(clk), .RN(n3758), .Q(
        \CACHE[1][136] ), .QN(n863) );
  DFFRX1 \CACHE_reg[1][135]  ( .D(n2102), .CK(clk), .RN(n3758), .Q(
        \CACHE[1][135] ), .QN(n862) );
  DFFRX1 \CACHE_reg[1][134]  ( .D(n2101), .CK(clk), .RN(n3758), .QN(n861) );
  DFFRX1 \CACHE_reg[1][133]  ( .D(n2100), .CK(clk), .RN(n3758), .QN(n860) );
  DFFRX1 \CACHE_reg[1][132]  ( .D(n2099), .CK(clk), .RN(n3757), .Q(
        \CACHE[1][132] ), .QN(n859) );
  DFFRX1 \CACHE_reg[1][131]  ( .D(n2098), .CK(clk), .RN(n3757), .Q(
        \CACHE[1][131] ), .QN(n858) );
  DFFRX1 \CACHE_reg[1][130]  ( .D(n2097), .CK(clk), .RN(n3757), .QN(n857) );
  DFFRX1 \CACHE_reg[1][129]  ( .D(n2096), .CK(clk), .RN(n3757), .Q(
        \CACHE[1][129] ), .QN(n856) );
  DFFRX1 \CACHE_reg[1][128]  ( .D(n2095), .CK(clk), .RN(n3757), .Q(
        \CACHE[1][128] ), .QN(n855) );
  DFFRX1 \CACHE_reg[4][154]  ( .D(n2586), .CK(clk), .RN(n3798), .QN(n1346) );
  DFFRX1 \CACHE_reg[4][153]  ( .D(n2585), .CK(clk), .RN(n3798), .Q(
        \CACHE[4][153] ), .QN(n1345) );
  DFFRX1 \CACHE_reg[4][152]  ( .D(n2584), .CK(clk), .RN(n3798), .QN(n1344) );
  DFFRX1 \CACHE_reg[4][151]  ( .D(n2583), .CK(clk), .RN(n3798), .QN(n1343) );
  DFFRX1 \CACHE_reg[4][150]  ( .D(n2582), .CK(clk), .RN(n3798), .QN(n1342) );
  DFFRX1 \CACHE_reg[4][149]  ( .D(n2581), .CK(clk), .RN(n3798), .Q(
        \CACHE[4][149] ), .QN(n1341) );
  DFFRX1 \CACHE_reg[4][148]  ( .D(n2580), .CK(clk), .RN(n3798), .Q(
        \CACHE[4][148] ), .QN(n1340) );
  DFFRX1 \CACHE_reg[4][147]  ( .D(n2579), .CK(clk), .RN(n3797), .QN(n1339) );
  DFFRX1 \CACHE_reg[4][146]  ( .D(n2578), .CK(clk), .RN(n3797), .QN(n1338) );
  DFFRX1 \CACHE_reg[4][145]  ( .D(n2577), .CK(clk), .RN(n3797), .QN(n1337) );
  DFFRX1 \CACHE_reg[4][144]  ( .D(n2576), .CK(clk), .RN(n3797), .QN(n1336) );
  DFFRX1 \CACHE_reg[4][143]  ( .D(n2575), .CK(clk), .RN(n3797), .Q(
        \CACHE[4][143] ), .QN(n1335) );
  DFFRX1 \CACHE_reg[4][142]  ( .D(n2574), .CK(clk), .RN(n3797), .Q(
        \CACHE[4][142] ), .QN(n1334) );
  DFFRX1 \CACHE_reg[4][141]  ( .D(n2573), .CK(clk), .RN(n3797), .Q(
        \CACHE[4][141] ), .QN(n1333) );
  DFFRX1 \CACHE_reg[4][140]  ( .D(n2572), .CK(clk), .RN(n3797), .QN(n1332) );
  DFFRX1 \CACHE_reg[4][139]  ( .D(n2571), .CK(clk), .RN(n3797), .Q(
        \CACHE[4][139] ), .QN(n1331) );
  DFFRX1 \CACHE_reg[4][138]  ( .D(n2570), .CK(clk), .RN(n3797), .Q(
        \CACHE[4][138] ), .QN(n1330) );
  DFFRX1 \CACHE_reg[4][137]  ( .D(n2569), .CK(clk), .RN(n3797), .Q(
        \CACHE[4][137] ), .QN(n1329) );
  DFFRX1 \CACHE_reg[4][136]  ( .D(n2568), .CK(clk), .RN(n3797), .Q(
        \CACHE[4][136] ), .QN(n1328) );
  DFFRX1 \CACHE_reg[4][135]  ( .D(n2567), .CK(clk), .RN(n3796), .QN(n1327) );
  DFFRX1 \CACHE_reg[4][134]  ( .D(n2566), .CK(clk), .RN(n3796), .QN(n1326) );
  DFFRX1 \CACHE_reg[4][133]  ( .D(n2565), .CK(clk), .RN(n3796), .QN(n1325) );
  DFFRX1 \CACHE_reg[4][132]  ( .D(n2564), .CK(clk), .RN(n3796), .Q(
        \CACHE[4][132] ), .QN(n1324) );
  DFFRX1 \CACHE_reg[4][131]  ( .D(n2563), .CK(clk), .RN(n3796), .Q(
        \CACHE[4][131] ), .QN(n1323) );
  DFFRX1 \CACHE_reg[4][130]  ( .D(n2562), .CK(clk), .RN(n3796), .QN(n1322) );
  DFFRX1 \CACHE_reg[4][129]  ( .D(n2561), .CK(clk), .RN(n3796), .Q(
        \CACHE[4][129] ), .QN(n1321) );
  DFFRX1 \CACHE_reg[4][128]  ( .D(n2560), .CK(clk), .RN(n3796), .Q(
        \CACHE[4][128] ), .QN(n1320) );
  DFFRX1 \CACHE_reg[0][154]  ( .D(n1966), .CK(clk), .RN(n3746), .QN(n726) );
  DFFRX1 \CACHE_reg[0][153]  ( .D(n1965), .CK(clk), .RN(n3746), .Q(
        \CACHE[0][153] ), .QN(n725) );
  DFFRX1 \CACHE_reg[0][152]  ( .D(n1964), .CK(clk), .RN(n3746), .QN(n724) );
  DFFRX1 \CACHE_reg[0][151]  ( .D(n1963), .CK(clk), .RN(n3746), .QN(n723) );
  DFFRX1 \CACHE_reg[0][150]  ( .D(n1962), .CK(clk), .RN(n3746), .QN(n722) );
  DFFRX1 \CACHE_reg[0][149]  ( .D(n1961), .CK(clk), .RN(n3746), .Q(
        \CACHE[0][149] ), .QN(n721) );
  DFFRX1 \CACHE_reg[0][148]  ( .D(n1960), .CK(clk), .RN(n3746), .Q(
        \CACHE[0][148] ), .QN(n720) );
  DFFRX1 \CACHE_reg[0][147]  ( .D(n1959), .CK(clk), .RN(n3746), .QN(n719) );
  DFFRX1 \CACHE_reg[0][146]  ( .D(n1958), .CK(clk), .RN(n3746), .QN(n718) );
  DFFRX1 \CACHE_reg[0][145]  ( .D(n1957), .CK(clk), .RN(n3746), .QN(n717) );
  DFFRX1 \CACHE_reg[0][144]  ( .D(n1956), .CK(clk), .RN(n3746), .QN(n716) );
  DFFRX1 \CACHE_reg[0][143]  ( .D(n1955), .CK(clk), .RN(n3745), .Q(
        \CACHE[0][143] ), .QN(n715) );
  DFFRX1 \CACHE_reg[0][142]  ( .D(n1954), .CK(clk), .RN(n3745), .Q(
        \CACHE[0][142] ), .QN(n714) );
  DFFRX1 \CACHE_reg[0][141]  ( .D(n1953), .CK(clk), .RN(n3745), .Q(
        \CACHE[0][141] ), .QN(n713) );
  DFFRX1 \CACHE_reg[0][140]  ( .D(n1952), .CK(clk), .RN(n3745), .QN(n712) );
  DFFRX1 \CACHE_reg[0][139]  ( .D(n1951), .CK(clk), .RN(n3745), .Q(
        \CACHE[0][139] ), .QN(n711) );
  DFFRX1 \CACHE_reg[0][138]  ( .D(n1950), .CK(clk), .RN(n3745), .Q(
        \CACHE[0][138] ), .QN(n710) );
  DFFRX1 \CACHE_reg[0][137]  ( .D(n1949), .CK(clk), .RN(n3745), .Q(
        \CACHE[0][137] ), .QN(n709) );
  DFFRX1 \CACHE_reg[0][136]  ( .D(n1948), .CK(clk), .RN(n3745), .Q(
        \CACHE[0][136] ), .QN(n708) );
  DFFRX1 \CACHE_reg[0][135]  ( .D(n1947), .CK(clk), .RN(n3745), .Q(
        \CACHE[0][135] ), .QN(n707) );
  DFFRX1 \CACHE_reg[0][134]  ( .D(n1946), .CK(clk), .RN(n3745), .QN(n706) );
  DFFRX1 \CACHE_reg[0][133]  ( .D(n1945), .CK(clk), .RN(n3745), .QN(n705) );
  DFFRX1 \CACHE_reg[0][132]  ( .D(n1944), .CK(clk), .RN(n3745), .Q(
        \CACHE[0][132] ), .QN(n704) );
  DFFRX1 \CACHE_reg[0][131]  ( .D(n1943), .CK(clk), .RN(n3744), .Q(
        \CACHE[0][131] ), .QN(n703) );
  DFFRX1 \CACHE_reg[0][130]  ( .D(n1942), .CK(clk), .RN(n3744), .QN(n702) );
  DFFRX1 \CACHE_reg[0][129]  ( .D(n1941), .CK(clk), .RN(n3744), .Q(
        \CACHE[0][129] ), .QN(n701) );
  DFFRX1 \CACHE_reg[0][128]  ( .D(n1940), .CK(clk), .RN(n3744), .Q(
        \CACHE[0][128] ), .QN(n700) );
  DFFRX1 \CACHE_reg[6][154]  ( .D(n2896), .CK(clk), .RN(n3824), .QN(n1656) );
  DFFRX1 \CACHE_reg[6][153]  ( .D(n2895), .CK(clk), .RN(n3824), .Q(
        \CACHE[6][153] ), .QN(n1655) );
  DFFRX1 \CACHE_reg[6][152]  ( .D(n2894), .CK(clk), .RN(n3824), .QN(n1654) );
  DFFRX1 \CACHE_reg[6][151]  ( .D(n2893), .CK(clk), .RN(n3824), .QN(n1653) );
  DFFRX1 \CACHE_reg[6][150]  ( .D(n2892), .CK(clk), .RN(n3824), .QN(n1652) );
  DFFRX1 \CACHE_reg[6][149]  ( .D(n2891), .CK(clk), .RN(n3823), .Q(
        \CACHE[6][149] ), .QN(n1651) );
  DFFRX1 \CACHE_reg[6][148]  ( .D(n2890), .CK(clk), .RN(n3823), .Q(
        \CACHE[6][148] ), .QN(n1650) );
  DFFRX1 \CACHE_reg[6][147]  ( .D(n2889), .CK(clk), .RN(n3823), .QN(n1649) );
  DFFRX1 \CACHE_reg[6][146]  ( .D(n2888), .CK(clk), .RN(n3823), .QN(n1648) );
  DFFRX1 \CACHE_reg[6][145]  ( .D(n2887), .CK(clk), .RN(n3823), .QN(n1647) );
  DFFRX1 \CACHE_reg[6][144]  ( .D(n2886), .CK(clk), .RN(n3823), .QN(n1646) );
  DFFRX1 \CACHE_reg[6][143]  ( .D(n2885), .CK(clk), .RN(n3823), .Q(
        \CACHE[6][143] ), .QN(n1645) );
  DFFRX1 \CACHE_reg[6][142]  ( .D(n2884), .CK(clk), .RN(n3823), .Q(
        \CACHE[6][142] ), .QN(n1644) );
  DFFRX1 \CACHE_reg[6][141]  ( .D(n2883), .CK(clk), .RN(n3823), .Q(
        \CACHE[6][141] ), .QN(n1643) );
  DFFRX1 \CACHE_reg[6][140]  ( .D(n2882), .CK(clk), .RN(n3823), .QN(n1642) );
  DFFRX1 \CACHE_reg[6][139]  ( .D(n2881), .CK(clk), .RN(n3823), .Q(
        \CACHE[6][139] ), .QN(n1641) );
  DFFRX1 \CACHE_reg[6][138]  ( .D(n2880), .CK(clk), .RN(n3823), .Q(
        \CACHE[6][138] ), .QN(n1640) );
  DFFRX1 \CACHE_reg[6][137]  ( .D(n2879), .CK(clk), .RN(n3822), .Q(
        \CACHE[6][137] ), .QN(n1639) );
  DFFRX1 \CACHE_reg[6][136]  ( .D(n2878), .CK(clk), .RN(n3822), .Q(
        \CACHE[6][136] ), .QN(n1638) );
  DFFRX1 \CACHE_reg[6][135]  ( .D(n2877), .CK(clk), .RN(n3822), .QN(n1637) );
  DFFRX1 \CACHE_reg[6][134]  ( .D(n2876), .CK(clk), .RN(n3822), .QN(n1636) );
  DFFRX1 \CACHE_reg[6][133]  ( .D(n2875), .CK(clk), .RN(n3822), .QN(n1635) );
  DFFRX1 \CACHE_reg[6][132]  ( .D(n2874), .CK(clk), .RN(n3822), .Q(
        \CACHE[6][132] ), .QN(n1634) );
  DFFRX1 \CACHE_reg[6][131]  ( .D(n2873), .CK(clk), .RN(n3822), .Q(
        \CACHE[6][131] ), .QN(n1633) );
  DFFRX1 \CACHE_reg[6][130]  ( .D(n2872), .CK(clk), .RN(n3822), .QN(n1632) );
  DFFRX1 \CACHE_reg[6][129]  ( .D(n2871), .CK(clk), .RN(n3822), .Q(
        \CACHE[6][129] ), .QN(n1631) );
  DFFRX1 \CACHE_reg[6][128]  ( .D(n2870), .CK(clk), .RN(n3822), .Q(
        \CACHE[6][128] ), .QN(n1630) );
  DFFRX1 \CACHE_reg[2][154]  ( .D(n2276), .CK(clk), .RN(n3772), .QN(n1036) );
  DFFRX1 \CACHE_reg[2][153]  ( .D(n2275), .CK(clk), .RN(n3772), .Q(
        \CACHE[2][153] ), .QN(n1035) );
  DFFRX1 \CACHE_reg[2][152]  ( .D(n2274), .CK(clk), .RN(n3772), .QN(n1034) );
  DFFRX1 \CACHE_reg[2][151]  ( .D(n2273), .CK(clk), .RN(n3772), .QN(n1033) );
  DFFRX1 \CACHE_reg[2][150]  ( .D(n2272), .CK(clk), .RN(n3772), .QN(n1032) );
  DFFRX1 \CACHE_reg[2][149]  ( .D(n2271), .CK(clk), .RN(n3772), .Q(
        \CACHE[2][149] ), .QN(n1031) );
  DFFRX1 \CACHE_reg[2][148]  ( .D(n2270), .CK(clk), .RN(n3772), .Q(
        \CACHE[2][148] ), .QN(n1030) );
  DFFRX1 \CACHE_reg[2][147]  ( .D(n2269), .CK(clk), .RN(n3772), .QN(n1029) );
  DFFRX1 \CACHE_reg[2][146]  ( .D(n2268), .CK(clk), .RN(n3772), .QN(n1028) );
  DFFRX1 \CACHE_reg[2][145]  ( .D(n2267), .CK(clk), .RN(n3771), .QN(n1027) );
  DFFRX1 \CACHE_reg[2][144]  ( .D(n2266), .CK(clk), .RN(n3771), .QN(n1026) );
  DFFRX1 \CACHE_reg[2][143]  ( .D(n2265), .CK(clk), .RN(n3771), .Q(
        \CACHE[2][143] ), .QN(n1025) );
  DFFRX1 \CACHE_reg[2][142]  ( .D(n2264), .CK(clk), .RN(n3771), .Q(
        \CACHE[2][142] ), .QN(n1024) );
  DFFRX1 \CACHE_reg[2][141]  ( .D(n2263), .CK(clk), .RN(n3771), .Q(
        \CACHE[2][141] ), .QN(n1023) );
  DFFRX1 \CACHE_reg[2][140]  ( .D(n2262), .CK(clk), .RN(n3771), .QN(n1022) );
  DFFRX1 \CACHE_reg[2][139]  ( .D(n2261), .CK(clk), .RN(n3771), .Q(
        \CACHE[2][139] ), .QN(n1021) );
  DFFRX1 \CACHE_reg[2][138]  ( .D(n2260), .CK(clk), .RN(n3771), .Q(
        \CACHE[2][138] ), .QN(n1020) );
  DFFRX1 \CACHE_reg[2][137]  ( .D(n2259), .CK(clk), .RN(n3771), .Q(
        \CACHE[2][137] ), .QN(n1019) );
  DFFRX1 \CACHE_reg[2][136]  ( .D(n2258), .CK(clk), .RN(n3771), .Q(
        \CACHE[2][136] ), .QN(n1018) );
  DFFRX1 \CACHE_reg[2][135]  ( .D(n2257), .CK(clk), .RN(n3771), .Q(
        \CACHE[2][135] ), .QN(n1017) );
  DFFRX1 \CACHE_reg[2][134]  ( .D(n2256), .CK(clk), .RN(n3771), .QN(n1016) );
  DFFRX1 \CACHE_reg[2][133]  ( .D(n2255), .CK(clk), .RN(n3770), .QN(n1015) );
  DFFRX1 \CACHE_reg[2][132]  ( .D(n2254), .CK(clk), .RN(n3770), .Q(
        \CACHE[2][132] ), .QN(n1014) );
  DFFRX1 \CACHE_reg[2][131]  ( .D(n2253), .CK(clk), .RN(n3770), .Q(
        \CACHE[2][131] ), .QN(n1013) );
  DFFRX1 \CACHE_reg[2][130]  ( .D(n2252), .CK(clk), .RN(n3770), .QN(n1012) );
  DFFRX1 \CACHE_reg[2][129]  ( .D(n2251), .CK(clk), .RN(n3770), .Q(
        \CACHE[2][129] ), .QN(n1011) );
  DFFRX1 \CACHE_reg[2][128]  ( .D(n2250), .CK(clk), .RN(n3770), .Q(
        \CACHE[2][128] ), .QN(n1010) );
  DFFRX1 \CACHE_reg[6][127]  ( .D(n2869), .CK(clk), .RN(n3822), .Q(
        \CACHE[6][127] ), .QN(n1629) );
  DFFRX1 \CACHE_reg[2][127]  ( .D(n2249), .CK(clk), .RN(n3770), .Q(
        \CACHE[2][127] ), .QN(n1009) );
  DFFRX1 \CACHE_reg[5][127]  ( .D(n2714), .CK(clk), .RN(n3809), .Q(
        \CACHE[5][127] ), .QN(n1474) );
  DFFRX1 \CACHE_reg[1][127]  ( .D(n2094), .CK(clk), .RN(n3757), .Q(
        \CACHE[1][127] ), .QN(n854) );
  DFFRX1 \CACHE_reg[7][127]  ( .D(n3024), .CK(clk), .RN(n3835), .Q(
        \CACHE[7][127] ), .QN(n1784) );
  DFFRX1 \CACHE_reg[3][127]  ( .D(n2404), .CK(clk), .RN(n3783), .Q(
        \CACHE[3][127] ), .QN(n1164) );
  DFFRX1 \CACHE_reg[4][127]  ( .D(n2559), .CK(clk), .RN(n3796), .Q(
        \CACHE[4][127] ), .QN(n1319) );
  DFFRX1 \CACHE_reg[0][127]  ( .D(n1939), .CK(clk), .RN(n3744), .Q(
        \CACHE[0][127] ), .QN(n699) );
  DFFRX1 \CACHE_reg[6][126]  ( .D(n2868), .CK(clk), .RN(n3822), .Q(
        \CACHE[6][126] ), .QN(n1628) );
  DFFRX1 \CACHE_reg[6][125]  ( .D(n2867), .CK(clk), .RN(n3821), .Q(
        \CACHE[6][125] ), .QN(n1627) );
  DFFRX1 \CACHE_reg[6][124]  ( .D(n2866), .CK(clk), .RN(n3821), .Q(
        \CACHE[6][124] ), .QN(n1626) );
  DFFRX1 \CACHE_reg[6][123]  ( .D(n2865), .CK(clk), .RN(n3821), .Q(
        \CACHE[6][123] ), .QN(n1625) );
  DFFRX1 \CACHE_reg[2][126]  ( .D(n2248), .CK(clk), .RN(n3770), .Q(
        \CACHE[2][126] ), .QN(n1008) );
  DFFRX1 \CACHE_reg[2][125]  ( .D(n2247), .CK(clk), .RN(n3770), .Q(
        \CACHE[2][125] ), .QN(n1007) );
  DFFRX1 \CACHE_reg[2][124]  ( .D(n2246), .CK(clk), .RN(n3770), .Q(
        \CACHE[2][124] ), .QN(n1006) );
  DFFRX1 \CACHE_reg[2][123]  ( .D(n2245), .CK(clk), .RN(n3770), .Q(
        \CACHE[2][123] ), .QN(n1005) );
  DFFRX1 \CACHE_reg[2][122]  ( .D(n2244), .CK(clk), .RN(n3770), .Q(
        \CACHE[2][122] ), .QN(n1004) );
  DFFRX1 \CACHE_reg[5][126]  ( .D(n2713), .CK(clk), .RN(n3809), .Q(
        \CACHE[5][126] ), .QN(n1473) );
  DFFRX1 \CACHE_reg[5][125]  ( .D(n2712), .CK(clk), .RN(n3809), .Q(
        \CACHE[5][125] ), .QN(n1472) );
  DFFRX1 \CACHE_reg[5][124]  ( .D(n2711), .CK(clk), .RN(n3808), .Q(
        \CACHE[5][124] ), .QN(n1471) );
  DFFRX1 \CACHE_reg[5][123]  ( .D(n2710), .CK(clk), .RN(n3808), .Q(
        \CACHE[5][123] ), .QN(n1470) );
  DFFRX1 \CACHE_reg[1][126]  ( .D(n2093), .CK(clk), .RN(n3757), .Q(
        \CACHE[1][126] ), .QN(n853) );
  DFFRX1 \CACHE_reg[1][125]  ( .D(n2092), .CK(clk), .RN(n3757), .Q(
        \CACHE[1][125] ), .QN(n852) );
  DFFRX1 \CACHE_reg[1][124]  ( .D(n2091), .CK(clk), .RN(n3757), .Q(
        \CACHE[1][124] ), .QN(n851) );
  DFFRX1 \CACHE_reg[1][123]  ( .D(n2090), .CK(clk), .RN(n3757), .Q(
        \CACHE[1][123] ), .QN(n850) );
  DFFRX1 \CACHE_reg[1][122]  ( .D(n2089), .CK(clk), .RN(n3757), .Q(
        \CACHE[1][122] ), .QN(n849) );
  DFFRX1 \CACHE_reg[7][126]  ( .D(n3023), .CK(clk), .RN(n3834), .Q(
        \CACHE[7][126] ), .QN(n1783) );
  DFFRX1 \CACHE_reg[7][125]  ( .D(n3022), .CK(clk), .RN(n3834), .Q(
        \CACHE[7][125] ), .QN(n1782) );
  DFFRX1 \CACHE_reg[7][124]  ( .D(n3021), .CK(clk), .RN(n3834), .Q(
        \CACHE[7][124] ), .QN(n1781) );
  DFFRX1 \CACHE_reg[7][123]  ( .D(n3020), .CK(clk), .RN(n3834), .Q(
        \CACHE[7][123] ), .QN(n1780) );
  DFFRX1 \CACHE_reg[3][126]  ( .D(n2403), .CK(clk), .RN(n3783), .Q(
        \CACHE[3][126] ), .QN(n1163) );
  DFFRX1 \CACHE_reg[3][125]  ( .D(n2402), .CK(clk), .RN(n3783), .Q(
        \CACHE[3][125] ), .QN(n1162) );
  DFFRX1 \CACHE_reg[3][124]  ( .D(n2401), .CK(clk), .RN(n3783), .Q(
        \CACHE[3][124] ), .QN(n1161) );
  DFFRX1 \CACHE_reg[3][123]  ( .D(n2400), .CK(clk), .RN(n3783), .Q(
        \CACHE[3][123] ), .QN(n1160) );
  DFFRX1 \CACHE_reg[3][122]  ( .D(n2399), .CK(clk), .RN(n3782), .Q(
        \CACHE[3][122] ), .QN(n1159) );
  DFFRX1 \CACHE_reg[4][126]  ( .D(n2558), .CK(clk), .RN(n3796), .Q(
        \CACHE[4][126] ), .QN(n1318) );
  DFFRX1 \CACHE_reg[4][125]  ( .D(n2557), .CK(clk), .RN(n3796), .Q(
        \CACHE[4][125] ), .QN(n1317) );
  DFFRX1 \CACHE_reg[4][124]  ( .D(n2556), .CK(clk), .RN(n3796), .Q(
        \CACHE[4][124] ), .QN(n1316) );
  DFFRX1 \CACHE_reg[4][123]  ( .D(n2555), .CK(clk), .RN(n3795), .Q(
        \CACHE[4][123] ), .QN(n1315) );
  DFFRX1 \CACHE_reg[0][126]  ( .D(n1938), .CK(clk), .RN(n3744), .Q(
        \CACHE[0][126] ), .QN(n698) );
  DFFRX1 \CACHE_reg[0][125]  ( .D(n1937), .CK(clk), .RN(n3744), .Q(
        \CACHE[0][125] ), .QN(n697) );
  DFFRX1 \CACHE_reg[0][124]  ( .D(n1936), .CK(clk), .RN(n3744), .Q(
        \CACHE[0][124] ), .QN(n696) );
  DFFRX1 \CACHE_reg[0][123]  ( .D(n1935), .CK(clk), .RN(n3744), .Q(
        \CACHE[0][123] ), .QN(n695) );
  DFFRX1 \CACHE_reg[0][122]  ( .D(n1934), .CK(clk), .RN(n3744), .Q(
        \CACHE[0][122] ), .QN(n694) );
  DFFRX1 \CACHE_reg[5][122]  ( .D(n2709), .CK(clk), .RN(n3808), .Q(
        \CACHE[5][122] ), .QN(n1469) );
  DFFRX1 \CACHE_reg[5][121]  ( .D(n2708), .CK(clk), .RN(n3808), .Q(
        \CACHE[5][121] ), .QN(n1468) );
  DFFRX1 \CACHE_reg[5][120]  ( .D(n2707), .CK(clk), .RN(n3808), .Q(
        \CACHE[5][120] ), .QN(n1467) );
  DFFRX1 \CACHE_reg[5][119]  ( .D(n2706), .CK(clk), .RN(n3808), .Q(
        \CACHE[5][119] ), .QN(n1466) );
  DFFRX1 \CACHE_reg[1][121]  ( .D(n2088), .CK(clk), .RN(n3757), .Q(
        \CACHE[1][121] ), .QN(n848) );
  DFFRX1 \CACHE_reg[1][120]  ( .D(n2087), .CK(clk), .RN(n3756), .Q(
        \CACHE[1][120] ), .QN(n847) );
  DFFRX1 \CACHE_reg[1][119]  ( .D(n2086), .CK(clk), .RN(n3756), .Q(
        \CACHE[1][119] ), .QN(n846) );
  DFFRX1 \CACHE_reg[6][122]  ( .D(n2864), .CK(clk), .RN(n3821), .Q(
        \CACHE[6][122] ), .QN(n1624) );
  DFFRX1 \CACHE_reg[6][121]  ( .D(n2863), .CK(clk), .RN(n3821), .Q(
        \CACHE[6][121] ), .QN(n1623) );
  DFFRX1 \CACHE_reg[6][120]  ( .D(n2862), .CK(clk), .RN(n3821), .Q(
        \CACHE[6][120] ), .QN(n1622) );
  DFFRX1 \CACHE_reg[6][119]  ( .D(n2861), .CK(clk), .RN(n3821), .Q(
        \CACHE[6][119] ), .QN(n1621) );
  DFFRX1 \CACHE_reg[2][121]  ( .D(n2243), .CK(clk), .RN(n3769), .Q(
        \CACHE[2][121] ), .QN(n1003) );
  DFFRX1 \CACHE_reg[2][120]  ( .D(n2242), .CK(clk), .RN(n3769), .Q(
        \CACHE[2][120] ), .QN(n1002) );
  DFFRX1 \CACHE_reg[2][119]  ( .D(n2241), .CK(clk), .RN(n3769), .Q(
        \CACHE[2][119] ), .QN(n1001) );
  DFFRX1 \CACHE_reg[4][122]  ( .D(n2554), .CK(clk), .RN(n3795), .Q(
        \CACHE[4][122] ), .QN(n1314) );
  DFFRX1 \CACHE_reg[4][121]  ( .D(n2553), .CK(clk), .RN(n3795), .Q(
        \CACHE[4][121] ), .QN(n1313) );
  DFFRX1 \CACHE_reg[4][120]  ( .D(n2552), .CK(clk), .RN(n3795), .Q(
        \CACHE[4][120] ), .QN(n1312) );
  DFFRX1 \CACHE_reg[4][119]  ( .D(n2551), .CK(clk), .RN(n3795), .Q(
        \CACHE[4][119] ), .QN(n1311) );
  DFFRX1 \CACHE_reg[0][121]  ( .D(n1933), .CK(clk), .RN(n3744), .Q(
        \CACHE[0][121] ), .QN(n693) );
  DFFRX1 \CACHE_reg[0][120]  ( .D(n1932), .CK(clk), .RN(n3744), .Q(
        \CACHE[0][120] ), .QN(n692) );
  DFFRX1 \CACHE_reg[0][119]  ( .D(n1931), .CK(clk), .RN(n3743), .Q(
        \CACHE[0][119] ), .QN(n691) );
  DFFRX1 \CACHE_reg[7][122]  ( .D(n3019), .CK(clk), .RN(n3834), .Q(
        \CACHE[7][122] ), .QN(n1779) );
  DFFRX1 \CACHE_reg[7][121]  ( .D(n3018), .CK(clk), .RN(n3834), .Q(
        \CACHE[7][121] ), .QN(n1778) );
  DFFRX1 \CACHE_reg[7][120]  ( .D(n3017), .CK(clk), .RN(n3834), .Q(
        \CACHE[7][120] ), .QN(n1777) );
  DFFRX1 \CACHE_reg[7][119]  ( .D(n3016), .CK(clk), .RN(n3834), .Q(
        \CACHE[7][119] ), .QN(n1776) );
  DFFRX1 \CACHE_reg[3][121]  ( .D(n2398), .CK(clk), .RN(n3782), .Q(
        \CACHE[3][121] ), .QN(n1158) );
  DFFRX1 \CACHE_reg[3][120]  ( .D(n2397), .CK(clk), .RN(n3782), .Q(
        \CACHE[3][120] ), .QN(n1157) );
  DFFRX1 \CACHE_reg[3][119]  ( .D(n2396), .CK(clk), .RN(n3782), .Q(
        \CACHE[3][119] ), .QN(n1156) );
  DFFRX1 \CACHE_reg[0][36]  ( .D(n1848), .CK(clk), .RN(n4142), .Q(
        \CACHE[0][36] ), .QN(n608) );
  DFFRX1 \CACHE_reg[0][32]  ( .D(n1844), .CK(clk), .RN(n4142), .Q(
        \CACHE[0][32] ), .QN(n604) );
  DFFRX1 \CACHE_reg[2][1]  ( .D(n2123), .CK(clk), .RN(n4142), .Q(\CACHE[2][1] ), .QN(n883) );
  MXI4X1 U2000 ( .A(\CACHE[0][129] ), .B(\CACHE[1][129] ), .C(\CACHE[2][129] ), 
        .D(\CACHE[3][129] ), .S0(n3682), .S1(n3711), .Y(n3623) );
  INVX3 U2001 ( .A(N30), .Y(n4141) );
  BUFX8 U2002 ( .A(n241), .Y(n3053) );
  AOI21XL U2003 ( .A0(mem_rdata[31]), .A1(n3898), .B0(n428), .Y(n241) );
  CLKINVX4 U2004 ( .A(n240), .Y(n3054) );
  INVX4 U2005 ( .A(n3054), .Y(n3055) );
  INVX4 U2006 ( .A(n3054), .Y(n3056) );
  OAI22X1 U2007 ( .A0(n4166), .A1(n3880), .B0(n3266), .B1(n3878), .Y(n446) );
  BUFX2 U2008 ( .A(n433), .Y(n3880) );
  BUFX4 U2009 ( .A(n434), .Y(n3878) );
  CLKBUFX4 U2010 ( .A(n3882), .Y(n3884) );
  CLKINVX8 U2011 ( .A(n239), .Y(n3057) );
  INVX8 U2012 ( .A(n3057), .Y(n3058) );
  INVX8 U2013 ( .A(n3057), .Y(n3059) );
  CLKINVX8 U2014 ( .A(n238), .Y(n3060) );
  INVX8 U2015 ( .A(n3060), .Y(n3061) );
  INVX8 U2016 ( .A(n3060), .Y(n3062) );
  CLKINVX8 U2017 ( .A(n236), .Y(n3063) );
  INVX8 U2018 ( .A(n3063), .Y(n3064) );
  INVX8 U2019 ( .A(n3063), .Y(n3065) );
  CLKINVX8 U2020 ( .A(n235), .Y(n3066) );
  INVX8 U2021 ( .A(n3066), .Y(n3067) );
  INVX8 U2022 ( .A(n3066), .Y(n3068) );
  CLKINVX8 U2023 ( .A(n237), .Y(n3069) );
  INVX8 U2024 ( .A(n3069), .Y(n3070) );
  INVX8 U2025 ( .A(n3069), .Y(n3071) );
  CLKINVX8 U2026 ( .A(n234), .Y(n3072) );
  INVX8 U2027 ( .A(n3072), .Y(n3073) );
  INVX8 U2028 ( .A(n3072), .Y(n3074) );
  CLKBUFX8 U2029 ( .A(n355), .Y(n3075) );
  INVX4 U2030 ( .A(n3320), .Y(n229) );
  INVX4 U2031 ( .A(n3318), .Y(n223) );
  INVX4 U2032 ( .A(n3322), .Y(n222) );
  BUFX12 U2033 ( .A(n216), .Y(n3076) );
  BUFX12 U2034 ( .A(n215), .Y(n3077) );
  BUFX12 U2035 ( .A(n214), .Y(n3078) );
  BUFX12 U2036 ( .A(n213), .Y(n3079) );
  BUFX12 U2037 ( .A(n209), .Y(n3080) );
  BUFX12 U2038 ( .A(n212), .Y(n3081) );
  BUFX12 U2039 ( .A(n221), .Y(n3082) );
  BUFX12 U2040 ( .A(n220), .Y(n3083) );
  BUFX12 U2041 ( .A(n219), .Y(n3084) );
  BUFX12 U2042 ( .A(n218), .Y(n3085) );
  BUFX12 U2043 ( .A(n217), .Y(n3086) );
  CLKBUFX8 U2044 ( .A(n468), .Y(n3087) );
  OAI22X1 U2045 ( .A0(n3892), .A1(n4152), .B0(n3363), .B1(n3075), .Y(n526) );
  OAI22X1 U2046 ( .A0(n4178), .A1(n3879), .B0(n3254), .B1(n3877), .Y(n432) );
  CLKBUFX4 U2047 ( .A(n433), .Y(n3879) );
  BUFX3 U2048 ( .A(n434), .Y(n3877) );
  BUFX12 U2049 ( .A(n273), .Y(n3088) );
  BUFX12 U2050 ( .A(n268), .Y(n3089) );
  BUFX12 U2051 ( .A(n302), .Y(n3090) );
  BUFX12 U2052 ( .A(n301), .Y(n3091) );
  BUFX12 U2053 ( .A(n300), .Y(n3092) );
  BUFX12 U2054 ( .A(n299), .Y(n3093) );
  BUFX12 U2055 ( .A(n305), .Y(n3094) );
  BUFX12 U2056 ( .A(n304), .Y(n3095) );
  BUFX12 U2057 ( .A(n303), .Y(n3096) );
  BUFX12 U2058 ( .A(n298), .Y(n3097) );
  BUFX12 U2059 ( .A(n272), .Y(n3098) );
  BUFX12 U2060 ( .A(n271), .Y(n3099) );
  BUFX12 U2061 ( .A(n270), .Y(n3100) );
  BUFX12 U2062 ( .A(n269), .Y(n3101) );
  BUFX12 U2063 ( .A(n267), .Y(n3102) );
  BUFX12 U2064 ( .A(n266), .Y(n3103) );
  BUFX12 U2065 ( .A(n265), .Y(n3104) );
  BUFX12 U2066 ( .A(n264), .Y(n3105) );
  BUFX12 U2067 ( .A(n263), .Y(n3106) );
  BUFX12 U2068 ( .A(n262), .Y(n3107) );
  BUFX12 U2069 ( .A(n261), .Y(n3108) );
  BUFX12 U2070 ( .A(n260), .Y(n3109) );
  BUFX12 U2071 ( .A(n259), .Y(n3110) );
  BUFX12 U2072 ( .A(n258), .Y(n3111) );
  BUFX12 U2073 ( .A(n257), .Y(n3112) );
  BUFX12 U2074 ( .A(n256), .Y(n3113) );
  BUFX12 U2075 ( .A(n255), .Y(n3114) );
  BUFX12 U2076 ( .A(n254), .Y(n3115) );
  BUFX12 U2077 ( .A(n253), .Y(n3116) );
  BUFX12 U2078 ( .A(n252), .Y(n3117) );
  BUFX12 U2079 ( .A(n251), .Y(n3118) );
  BUFX12 U2080 ( .A(n250), .Y(n3119) );
  BUFX12 U2081 ( .A(n249), .Y(n3120) );
  BUFX12 U2082 ( .A(n248), .Y(n3121) );
  BUFX12 U2083 ( .A(n247), .Y(n3122) );
  BUFX12 U2084 ( .A(n245), .Y(n3123) );
  BUFX12 U2085 ( .A(n244), .Y(n3124) );
  BUFX12 U2086 ( .A(n243), .Y(n3125) );
  BUFX12 U2087 ( .A(n228), .Y(n3126) );
  BUFX12 U2088 ( .A(n227), .Y(n3127) );
  BUFX12 U2089 ( .A(n226), .Y(n3128) );
  BUFX12 U2090 ( .A(n225), .Y(n3129) );
  BUFX12 U2091 ( .A(n224), .Y(n3130) );
  BUFX12 U2092 ( .A(n233), .Y(n3131) );
  BUFX12 U2093 ( .A(n232), .Y(n3132) );
  BUFX12 U2094 ( .A(n231), .Y(n3133) );
  BUFX12 U2095 ( .A(n230), .Y(n3134) );
  BUFX12 U2096 ( .A(n326), .Y(n3135) );
  BUFX12 U2097 ( .A(n324), .Y(n3136) );
  BUFX12 U2098 ( .A(n323), .Y(n3137) );
  BUFX12 U2099 ( .A(n322), .Y(n3138) );
  BUFX12 U2100 ( .A(n321), .Y(n3139) );
  BUFX12 U2101 ( .A(n327), .Y(n3140) );
  BUFX12 U2102 ( .A(n325), .Y(n3141) );
  BUFX12 U2103 ( .A(n320), .Y(n3142) );
  BUFX12 U2104 ( .A(n319), .Y(n3143) );
  BUFX12 U2105 ( .A(n318), .Y(n3144) );
  BUFX12 U2106 ( .A(n317), .Y(n3145) );
  BUFX12 U2107 ( .A(n316), .Y(n3146) );
  BUFX12 U2108 ( .A(n287), .Y(n3147) );
  BUFX12 U2109 ( .A(n286), .Y(n3148) );
  BUFX12 U2110 ( .A(n281), .Y(n3149) );
  BUFX12 U2111 ( .A(n279), .Y(n3150) );
  BUFX12 U2112 ( .A(n275), .Y(n3151) );
  BUFX12 U2113 ( .A(n274), .Y(n3152) );
  BUFX12 U2114 ( .A(n297), .Y(n3153) );
  BUFX12 U2115 ( .A(n296), .Y(n3154) );
  BUFX12 U2116 ( .A(n295), .Y(n3155) );
  BUFX12 U2117 ( .A(n291), .Y(n3156) );
  BUFX12 U2118 ( .A(n289), .Y(n3157) );
  BUFX12 U2119 ( .A(n288), .Y(n3158) );
  BUFX12 U2120 ( .A(n278), .Y(n3159) );
  BUFX12 U2121 ( .A(n292), .Y(n3160) );
  BUFX12 U2122 ( .A(n280), .Y(n3161) );
  BUFX12 U2123 ( .A(n293), .Y(n3162) );
  BUFX12 U2124 ( .A(n282), .Y(n3163) );
  BUFX12 U2125 ( .A(n294), .Y(n3164) );
  BUFX12 U2126 ( .A(n283), .Y(n3165) );
  BUFX12 U2127 ( .A(n290), .Y(n3166) );
  BUFX12 U2128 ( .A(n284), .Y(n3167) );
  BUFX12 U2129 ( .A(n276), .Y(n3168) );
  BUFX12 U2130 ( .A(n285), .Y(n3169) );
  BUFX12 U2131 ( .A(n277), .Y(n3170) );
  BUFX12 U2132 ( .A(n331), .Y(n3171) );
  BUFX12 U2133 ( .A(n328), .Y(n3172) );
  BUFX12 U2134 ( .A(n330), .Y(n3173) );
  BUFX12 U2135 ( .A(n178), .Y(n3174) );
  BUFX12 U2136 ( .A(n334), .Y(n3175) );
  BUFX12 U2137 ( .A(n309), .Y(n3176) );
  BUFX12 U2138 ( .A(n308), .Y(n3177) );
  BUFX12 U2139 ( .A(n307), .Y(n3178) );
  BUFX12 U2140 ( .A(n306), .Y(n3179) );
  BUFX12 U2141 ( .A(n329), .Y(n3180) );
  BUFX12 U2142 ( .A(n335), .Y(n3181) );
  BUFX12 U2143 ( .A(n315), .Y(n3182) );
  BUFX12 U2144 ( .A(n314), .Y(n3183) );
  BUFX12 U2145 ( .A(n313), .Y(n3184) );
  BUFX12 U2146 ( .A(n312), .Y(n3185) );
  BUFX12 U2147 ( .A(n311), .Y(n3186) );
  BUFX12 U2148 ( .A(n310), .Y(n3187) );
  BUFX12 U2149 ( .A(n333), .Y(n3188) );
  BUFX12 U2150 ( .A(n332), .Y(n3189) );
  NOR2X8 U2151 ( .A(n3336), .B(n356), .Y(n180) );
  NAND2X2 U2152 ( .A(n3337), .B(n3338), .Y(n356) );
  OAI31X4 U2153 ( .A0(n3341), .A1(n3315), .A2(n4146), .B0(n430), .Y(n434) );
  CLKINVX1 U2154 ( .A(n3342), .Y(n3341) );
  NAND2BX4 U2155 ( .AN(n429), .B(n361), .Y(n430) );
  OAI21X1 U2156 ( .A0(n3317), .A1(n4145), .B0(n3311), .Y(n532) );
  NOR2X2 U2157 ( .A(n363), .B(n533), .Y(n176) );
  INVX16 U2158 ( .A(n4139), .Y(n4138) );
  XNOR2X2 U2159 ( .A(N44), .B(proc_addr[20]), .Y(n564) );
  XNOR2X2 U2160 ( .A(N45), .B(proc_addr[19]), .Y(n563) );
  XNOR2X2 U2161 ( .A(N50), .B(proc_addr[14]), .Y(n562) );
  INVX3 U2162 ( .A(n429), .Y(n3342) );
  NAND3X1 U2163 ( .A(n3313), .B(n3314), .C(n4143), .Y(n433) );
  NAND3X1 U2164 ( .A(n3315), .B(n4146), .C(n4143), .Y(n467) );
  BUFX4 U2165 ( .A(n3718), .Y(n3689) );
  CLKBUFX3 U2166 ( .A(n3691), .Y(n3712) );
  NAND2X1 U2167 ( .A(N33), .B(n3317), .Y(n363) );
  CLKINVX1 U2168 ( .A(n3313), .Y(n4146) );
  NAND4X4 U2169 ( .A(n539), .B(n540), .C(n541), .D(n542), .Y(n533) );
  NOR4X2 U2170 ( .A(n543), .B(n544), .C(n545), .D(n546), .Y(n542) );
  NAND3X2 U2171 ( .A(n4144), .B(n3316), .C(proc_write), .Y(n361) );
  INVX12 U2172 ( .A(N31), .Y(n4139) );
  CLKMX2X2 U2173 ( .A(n3352), .B(n3353), .S0(n3726), .Y(N59) );
  MXI2X1 U2174 ( .A(n3623), .B(n3624), .S0(n3726), .Y(N58) );
  CLKMX2X2 U2175 ( .A(n3349), .B(n3350), .S0(n3727), .Y(N47) );
  CLKMX2X2 U2176 ( .A(n3347), .B(n3348), .S0(n3728), .Y(N43) );
  NAND2X1 U2177 ( .A(n3651), .B(n4137), .Y(n3381) );
  NAND2X1 U2178 ( .A(n3652), .B(n3728), .Y(n3382) );
  CLKMX2X2 U2179 ( .A(n3345), .B(n3346), .S0(n3728), .Y(N37) );
  MXI2X1 U2180 ( .A(n3655), .B(n3656), .S0(n3728), .Y(N35) );
  OAI22XL U2181 ( .A0(n3885), .A1(n4178), .B0(n3190), .B1(n3883), .Y(n365) );
  OAI2BB1X1 U2182 ( .A0N(mem_rdata[12]), .A1N(n3900), .B0(n3323), .Y(n3322) );
  OAI2BB1X1 U2183 ( .A0N(mem_rdata[13]), .A1N(n3900), .B0(n3319), .Y(n3318) );
  OAI2BB1X1 U2184 ( .A0N(mem_rdata[19]), .A1N(n3899), .B0(n3321), .Y(n3320) );
  NAND2X1 U2185 ( .A(n3324), .B(n3325), .Y(n2123) );
  NAND2X1 U2186 ( .A(n3328), .B(n3329), .Y(n1844) );
  NAND2X1 U2187 ( .A(n3326), .B(n3327), .Y(n1848) );
  BUFX4 U2188 ( .A(n3882), .Y(n3883) );
  INVX3 U2189 ( .A(N32), .Y(n4137) );
  INVX3 U2190 ( .A(n4137), .Y(n4136) );
  CLKBUFX3 U2191 ( .A(n3958), .Y(n3947) );
  NOR3X1 U2192 ( .A(n4138), .B(n4136), .C(n4140), .Y(n347) );
  NOR3X1 U2193 ( .A(n4139), .B(n4140), .C(n4137), .Y(n343) );
  NOR3X1 U2194 ( .A(n4140), .B(n4138), .C(n4137), .Y(n338) );
  NOR3X1 U2195 ( .A(n4140), .B(n4136), .C(n4139), .Y(n177) );
  BUFX4 U2196 ( .A(n368), .Y(n3882) );
  CLKMX2X2 U2197 ( .A(n3385), .B(n3386), .S0(n3723), .Y(n3190) );
  CLKMX2X2 U2198 ( .A(n3575), .B(n3576), .S0(n3719), .Y(n3191) );
  CLKMX2X2 U2199 ( .A(n3513), .B(n3514), .S0(n3723), .Y(n3192) );
  CLKMX2X2 U2200 ( .A(n3515), .B(n3516), .S0(n3723), .Y(n3193) );
  CLKMX2X2 U2201 ( .A(n3517), .B(n3518), .S0(n3723), .Y(n3194) );
  CLKMX2X2 U2202 ( .A(n3519), .B(n3520), .S0(n3723), .Y(n3195) );
  CLKMX2X2 U2203 ( .A(n3521), .B(n3522), .S0(n3723), .Y(n3196) );
  CLKMX2X2 U2204 ( .A(n3523), .B(n3524), .S0(n3723), .Y(n3197) );
  CLKMX2X2 U2205 ( .A(n3525), .B(n3526), .S0(n3723), .Y(n3198) );
  CLKMX2X2 U2206 ( .A(n3561), .B(n3562), .S0(n3725), .Y(n3199) );
  CLKMX2X2 U2207 ( .A(n3563), .B(n3564), .S0(n3725), .Y(n3200) );
  CLKMX2X2 U2208 ( .A(n3565), .B(n3566), .S0(n3725), .Y(n3201) );
  CLKMX2X2 U2209 ( .A(n3567), .B(n3568), .S0(n3725), .Y(n3202) );
  CLKMX2X2 U2210 ( .A(n3569), .B(n3570), .S0(n3725), .Y(n3203) );
  CLKMX2X2 U2211 ( .A(n3571), .B(n3572), .S0(n3725), .Y(n3204) );
  CLKMX2X2 U2212 ( .A(n3573), .B(n3574), .S0(n3725), .Y(n3205) );
  CLKMX2X2 U2213 ( .A(n3527), .B(n3528), .S0(n3724), .Y(n3206) );
  CLKMX2X2 U2214 ( .A(n3529), .B(n3530), .S0(n3724), .Y(n3207) );
  CLKMX2X2 U2215 ( .A(n3531), .B(n3532), .S0(n3724), .Y(n3208) );
  CLKMX2X2 U2216 ( .A(n3533), .B(n3534), .S0(n3724), .Y(n3209) );
  CLKMX2X2 U2217 ( .A(n3535), .B(n3536), .S0(n3724), .Y(n3210) );
  CLKMX2X2 U2218 ( .A(n3537), .B(n3538), .S0(n3724), .Y(n3211) );
  CLKMX2X2 U2219 ( .A(n3539), .B(n3540), .S0(n3724), .Y(n3212) );
  CLKMX2X2 U2220 ( .A(n3541), .B(n3542), .S0(n3724), .Y(n3213) );
  CLKMX2X2 U2221 ( .A(n3543), .B(n3544), .S0(n3724), .Y(n3214) );
  CLKMX2X2 U2222 ( .A(n3545), .B(n3546), .S0(n3724), .Y(n3215) );
  CLKMX2X2 U2223 ( .A(n3547), .B(n3548), .S0(n3724), .Y(n3216) );
  CLKMX2X2 U2224 ( .A(n3549), .B(n3550), .S0(n3724), .Y(n3217) );
  CLKMX2X2 U2225 ( .A(n3551), .B(n3552), .S0(n3725), .Y(n3218) );
  CLKMX2X2 U2226 ( .A(n3553), .B(n3554), .S0(n3725), .Y(n3219) );
  CLKMX2X2 U2227 ( .A(n3555), .B(n3556), .S0(n3725), .Y(n3220) );
  CLKMX2X2 U2228 ( .A(n3557), .B(n3558), .S0(n3725), .Y(n3221) );
  CLKMX2X2 U2229 ( .A(n3559), .B(n3560), .S0(n3725), .Y(n3222) );
  CLKMX2X2 U2230 ( .A(n3621), .B(n3622), .S0(n3726), .Y(n3223) );
  CLKMX2X2 U2231 ( .A(n3599), .B(n3600), .S0(n4136), .Y(n3224) );
  CLKMX2X2 U2232 ( .A(n3601), .B(n3602), .S0(n3724), .Y(n3225) );
  CLKMX2X2 U2233 ( .A(n3603), .B(n3604), .S0(n4136), .Y(n3226) );
  CLKMX2X2 U2234 ( .A(n3605), .B(n3606), .S0(n3724), .Y(n3227) );
  CLKMX2X2 U2235 ( .A(n3607), .B(n3608), .S0(n3720), .Y(n3228) );
  CLKMX2X2 U2236 ( .A(n3609), .B(n3610), .S0(n3721), .Y(n3229) );
  CLKMX2X2 U2237 ( .A(n3611), .B(n3612), .S0(n3719), .Y(n3230) );
  CLKMX2X2 U2238 ( .A(n3613), .B(n3614), .S0(n3719), .Y(n3231) );
  CLKMX2X2 U2239 ( .A(n3615), .B(n3616), .S0(n3719), .Y(n3232) );
  CLKMX2X2 U2240 ( .A(n3617), .B(n3618), .S0(n3728), .Y(n3233) );
  CLKMX2X2 U2241 ( .A(n3619), .B(n3620), .S0(n4136), .Y(n3234) );
  CLKMX2X2 U2242 ( .A(n3395), .B(n3396), .S0(n3720), .Y(n3235) );
  CLKMX2X2 U2243 ( .A(n3401), .B(n3402), .S0(n3722), .Y(n3236) );
  CLKMX2X2 U2244 ( .A(n3399), .B(n3400), .S0(n4136), .Y(n3237) );
  CLKMX2X2 U2245 ( .A(n3403), .B(n3404), .S0(n3723), .Y(n3238) );
  CLKMX2X2 U2246 ( .A(n3387), .B(n3388), .S0(n3725), .Y(n3239) );
  CLKMX2X2 U2247 ( .A(n3391), .B(n3392), .S0(n3724), .Y(n3240) );
  CLKMX2X2 U2248 ( .A(n3405), .B(n3406), .S0(n3724), .Y(n3241) );
  CLKMX2X2 U2249 ( .A(n3389), .B(n3390), .S0(n3719), .Y(n3242) );
  CLKMX2X2 U2250 ( .A(n3393), .B(n3394), .S0(n3719), .Y(n3243) );
  CLKMX2X2 U2251 ( .A(n3397), .B(n3398), .S0(n3721), .Y(n3244) );
  NOR3BXL U2252 ( .AN(n538), .B(n7), .C(n3311), .Y(n4179) );
  BUFX4 U2253 ( .A(n4179), .Y(mem_read) );
  AND2X2 U2254 ( .A(n3381), .B(n3382), .Y(n3245) );
  NAND2X1 U2255 ( .A(n3344), .B(n430), .Y(n368) );
  CLKMX2X2 U2256 ( .A(n3497), .B(n3498), .S0(n3722), .Y(n3246) );
  CLKMX2X2 U2257 ( .A(n3499), .B(n3500), .S0(n3722), .Y(n3247) );
  CLKMX2X2 U2258 ( .A(n3501), .B(n3502), .S0(n3722), .Y(n3248) );
  CLKMX2X2 U2259 ( .A(n3503), .B(n3504), .S0(n3723), .Y(n3249) );
  CLKMX2X2 U2260 ( .A(n3505), .B(n3506), .S0(n3723), .Y(n3250) );
  CLKMX2X2 U2261 ( .A(n3507), .B(n3508), .S0(n3723), .Y(n3251) );
  CLKMX2X2 U2262 ( .A(n3509), .B(n3510), .S0(n3723), .Y(n3252) );
  CLKMX2X2 U2263 ( .A(n3511), .B(n3512), .S0(n3723), .Y(n3253) );
  CLKMX2X2 U2264 ( .A(n3449), .B(n3450), .S0(n3722), .Y(n3254) );
  CLKMX2X2 U2265 ( .A(n3451), .B(n3452), .S0(n3725), .Y(n3255) );
  CLKMX2X2 U2266 ( .A(n3453), .B(n3454), .S0(n3722), .Y(n3256) );
  CLKMX2X2 U2267 ( .A(n3455), .B(n3456), .S0(n3721), .Y(n3257) );
  CLKMX2X2 U2268 ( .A(n3457), .B(n3458), .S0(n3721), .Y(n3258) );
  CLKMX2X2 U2269 ( .A(n3459), .B(n3460), .S0(n3721), .Y(n3259) );
  CLKMX2X2 U2270 ( .A(n3461), .B(n3462), .S0(n3721), .Y(n3260) );
  CLKMX2X2 U2271 ( .A(n3463), .B(n3464), .S0(n3721), .Y(n3261) );
  CLKMX2X2 U2272 ( .A(n3465), .B(n3466), .S0(n3721), .Y(n3262) );
  CLKMX2X2 U2273 ( .A(n3467), .B(n3468), .S0(n3721), .Y(n3263) );
  CLKMX2X2 U2274 ( .A(n3469), .B(n3470), .S0(n3721), .Y(n3264) );
  CLKMX2X2 U2275 ( .A(n3471), .B(n3472), .S0(n3721), .Y(n3265) );
  CLKMX2X2 U2276 ( .A(n3473), .B(n3474), .S0(n3721), .Y(n3266) );
  CLKMX2X2 U2277 ( .A(n3475), .B(n3476), .S0(n3721), .Y(n3267) );
  CLKMX2X2 U2278 ( .A(n3477), .B(n3478), .S0(n3721), .Y(n3268) );
  CLKMX2X2 U2279 ( .A(n3479), .B(n3480), .S0(n3722), .Y(n3269) );
  CLKMX2X2 U2280 ( .A(n3481), .B(n3482), .S0(n3722), .Y(n3270) );
  CLKMX2X2 U2281 ( .A(n3483), .B(n3484), .S0(n3722), .Y(n3271) );
  CLKMX2X2 U2282 ( .A(n3485), .B(n3486), .S0(n3722), .Y(n3272) );
  CLKMX2X2 U2283 ( .A(n3487), .B(n3488), .S0(n3722), .Y(n3273) );
  CLKMX2X2 U2284 ( .A(n3489), .B(n3490), .S0(n3722), .Y(n3274) );
  CLKMX2X2 U2285 ( .A(n3491), .B(n3492), .S0(n3722), .Y(n3275) );
  CLKMX2X2 U2286 ( .A(n3493), .B(n3494), .S0(n3722), .Y(n3276) );
  CLKMX2X2 U2287 ( .A(n3495), .B(n3496), .S0(n3722), .Y(n3277) );
  CLKMX2X2 U2288 ( .A(n3577), .B(n3578), .S0(N32), .Y(n3278) );
  CLKMX2X2 U2289 ( .A(n3579), .B(n3580), .S0(N32), .Y(n3279) );
  CLKMX2X2 U2290 ( .A(n3581), .B(n3582), .S0(N32), .Y(n3280) );
  CLKMX2X2 U2291 ( .A(n3583), .B(n3584), .S0(n4136), .Y(n3281) );
  CLKMX2X2 U2292 ( .A(n3585), .B(n3586), .S0(n4136), .Y(n3282) );
  CLKMX2X2 U2293 ( .A(n3587), .B(n3588), .S0(n4136), .Y(n3283) );
  CLKMX2X2 U2294 ( .A(n3589), .B(n3590), .S0(n4136), .Y(n3284) );
  CLKMX2X2 U2295 ( .A(n3591), .B(n3592), .S0(n4136), .Y(n3285) );
  CLKMX2X2 U2296 ( .A(n3593), .B(n3594), .S0(N32), .Y(n3286) );
  CLKMX2X2 U2297 ( .A(n3595), .B(n3596), .S0(N32), .Y(n3287) );
  CLKMX2X2 U2298 ( .A(n3597), .B(n3598), .S0(n4136), .Y(n3288) );
  CLKMX2X2 U2299 ( .A(n3433), .B(n3434), .S0(n3721), .Y(n3289) );
  CLKMX2X2 U2300 ( .A(n3435), .B(n3436), .S0(n3725), .Y(n3290) );
  CLKMX2X2 U2301 ( .A(n3437), .B(n3438), .S0(n3722), .Y(n3291) );
  CLKMX2X2 U2302 ( .A(n3439), .B(n3440), .S0(n3723), .Y(n3292) );
  CLKMX2X2 U2303 ( .A(n3441), .B(n3442), .S0(n3720), .Y(n3293) );
  CLKMX2X2 U2304 ( .A(n3443), .B(n3444), .S0(n3721), .Y(n3294) );
  CLKMX2X2 U2305 ( .A(n3445), .B(n3446), .S0(n3725), .Y(n3295) );
  CLKMX2X2 U2306 ( .A(n3447), .B(n3448), .S0(n3723), .Y(n3296) );
  CLKMX2X2 U2307 ( .A(n3407), .B(n3408), .S0(n3720), .Y(n3297) );
  CLKMX2X2 U2308 ( .A(n3413), .B(n3414), .S0(n3720), .Y(n3298) );
  CLKMX2X2 U2309 ( .A(n3415), .B(n3416), .S0(n3720), .Y(n3299) );
  CLKMX2X2 U2310 ( .A(n3417), .B(n3418), .S0(n3720), .Y(n3300) );
  CLKMX2X2 U2311 ( .A(n3419), .B(n3420), .S0(n3720), .Y(n3301) );
  CLKMX2X2 U2312 ( .A(n3421), .B(n3422), .S0(n3720), .Y(n3302) );
  CLKMX2X2 U2313 ( .A(n3425), .B(n3426), .S0(n3720), .Y(n3303) );
  CLKMX2X2 U2314 ( .A(n3427), .B(n3428), .S0(n3720), .Y(n3304) );
  CLKMX2X2 U2315 ( .A(n3429), .B(n3430), .S0(n3720), .Y(n3305) );
  CLKMX2X2 U2316 ( .A(n3431), .B(n3432), .S0(n3720), .Y(n3306) );
  CLKMX2X2 U2317 ( .A(n3409), .B(n3410), .S0(n3720), .Y(n3307) );
  CLKMX2X2 U2318 ( .A(n3411), .B(n3412), .S0(n3720), .Y(n3308) );
  CLKMX2X2 U2319 ( .A(n3423), .B(n3424), .S0(n3720), .Y(n3309) );
  CLKINVX1 U2320 ( .A(n535), .Y(n3873) );
  CLKBUFX3 U2321 ( .A(n3688), .Y(n3692) );
  CLKINVX1 U2322 ( .A(n3314), .Y(n3315) );
  CLKINVX1 U2323 ( .A(n3312), .Y(n3313) );
  CLKINVX1 U2324 ( .A(mem_ready), .Y(n3310) );
  INVX3 U2325 ( .A(n3310), .Y(n3311) );
  CLKINVX1 U2326 ( .A(proc_addr[0]), .Y(n3312) );
  CLKINVX1 U2327 ( .A(proc_addr[1]), .Y(n3314) );
  CLKINVX1 U2328 ( .A(proc_read), .Y(n3316) );
  INVX3 U2329 ( .A(n3316), .Y(n3317) );
  OA22XL U2330 ( .A0(n3886), .A1(n4165), .B0(n3308), .B1(n3884), .Y(n3319) );
  OA22XL U2331 ( .A0(n3886), .A1(n4159), .B0(n3309), .B1(n3884), .Y(n3321) );
  OA22XL U2332 ( .A0(n3886), .A1(n4166), .B0(n3307), .B1(n3884), .Y(n3323) );
  MXI2X2 U2333 ( .A(n3627), .B(n3628), .S0(n3727), .Y(N56) );
  MXI4XL U2334 ( .A(\CACHE[4][131] ), .B(\CACHE[5][131] ), .C(\CACHE[6][131] ), 
        .D(\CACHE[7][131] ), .S0(n3682), .S1(n3712), .Y(n3628) );
  MXI4XL U2335 ( .A(\CACHE[0][131] ), .B(\CACHE[1][131] ), .C(\CACHE[2][131] ), 
        .D(\CACHE[3][131] ), .S0(n3682), .S1(n3712), .Y(n3627) );
  CLKBUFX3 U2336 ( .A(n3690), .Y(n3714) );
  OR2X1 U2337 ( .A(n883), .B(n4101), .Y(n3324) );
  OR2XL U2338 ( .A(n211), .B(n4114), .Y(n3325) );
  AOI21X4 U2339 ( .A0(mem_rdata[1]), .A1(n3901), .B0(n369), .Y(n211) );
  BUFX2 U2340 ( .A(n4125), .Y(n4114) );
  BUFX20 U2341 ( .A(n3716), .Y(n3718) );
  OR2X1 U2342 ( .A(n608), .B(n3934), .Y(n3326) );
  OR2XL U2343 ( .A(n246), .B(n3947), .Y(n3327) );
  AOI21X4 U2344 ( .A0(mem_rdata[36]), .A1(n3898), .B0(n438), .Y(n246) );
  OR2X1 U2345 ( .A(n604), .B(n3933), .Y(n3328) );
  OR2XL U2346 ( .A(n242), .B(n3956), .Y(n3329) );
  AOI21X4 U2347 ( .A0(mem_rdata[32]), .A1(n3898), .B0(n432), .Y(n242) );
  CLKMX2X2 U2348 ( .A(n3330), .B(n3331), .S0(n3728), .Y(N36) );
  MXI4XL U2349 ( .A(n723), .B(n878), .C(n1033), .D(n1188), .S0(n3685), .S1(
        n3715), .Y(n3330) );
  MXI4XL U2350 ( .A(n1343), .B(n1498), .C(n1653), .D(n1808), .S0(n3685), .S1(
        n3715), .Y(n3331) );
  CLKMX2X2 U2351 ( .A(n3332), .B(n3333), .S0(n3728), .Y(N41) );
  MXI4XL U2352 ( .A(n718), .B(n873), .C(n1028), .D(n1183), .S0(n3684), .S1(
        n3714), .Y(n3332) );
  MXI4XL U2353 ( .A(n1338), .B(n1493), .C(n1648), .D(n1803), .S0(n3684), .S1(
        n3714), .Y(n3333) );
  CLKMX2X2 U2354 ( .A(n3334), .B(n3335), .S0(n3728), .Y(N40) );
  MXI4XL U2355 ( .A(n719), .B(n874), .C(n1029), .D(n1184), .S0(n3684), .S1(
        n3714), .Y(n3334) );
  MXI4XL U2356 ( .A(n1339), .B(n1494), .C(n1649), .D(n1804), .S0(n3684), .S1(
        n3714), .Y(n3335) );
  CLKBUFX2 U2357 ( .A(n3691), .Y(n3713) );
  CLKBUFX3 U2358 ( .A(n353), .Y(n3890) );
  BUFX20 U2359 ( .A(N30), .Y(n3660) );
  NAND3XL U2360 ( .A(n3342), .B(n3343), .C(n3312), .Y(n3344) );
  OAI22XL U2361 ( .A0(n699), .A1(n3941), .B0(n180), .B1(n3954), .Y(n1939) );
  OAI22XL U2362 ( .A0(n854), .A1(n3913), .B0(n180), .B1(n3927), .Y(n2094) );
  OAI22XL U2363 ( .A0(n1164), .A1(n4081), .B0(n180), .B1(n4095), .Y(n2404) );
  OAI22XL U2364 ( .A0(n1319), .A1(n4053), .B0(n180), .B1(n4066), .Y(n2559) );
  OAI22XL U2365 ( .A0(n1474), .A1(n4025), .B0(n180), .B1(n4039), .Y(n2714) );
  OAI22XL U2366 ( .A0(n1629), .A1(n3997), .B0(n180), .B1(n4010), .Y(n2869) );
  OAI22XL U2367 ( .A0(n1784), .A1(n3969), .B0(n180), .B1(n3983), .Y(n3024) );
  OAI22XL U2368 ( .A0(n1009), .A1(n4099), .B0(n180), .B1(n4113), .Y(n2249) );
  AND2X2 U2369 ( .A(mem_rdata[127]), .B(n3901), .Y(n3336) );
  OR2X1 U2370 ( .A(n3890), .B(n4147), .Y(n3337) );
  OR2XL U2371 ( .A(n3378), .B(n3075), .Y(n3338) );
  CLKMX2X2 U2372 ( .A(n3339), .B(n3340), .S0(n3728), .Y(N42) );
  MXI4XL U2373 ( .A(n717), .B(n872), .C(n1027), .D(n1182), .S0(n3684), .S1(
        n3714), .Y(n3339) );
  MXI4XL U2374 ( .A(n1337), .B(n1492), .C(n1647), .D(n1802), .S0(n3684), .S1(
        n3714), .Y(n3340) );
  BUFX8 U2375 ( .A(n3663), .Y(n3681) );
  AOI2BB2X1 U2376 ( .B0(n532), .B1(n533), .A0N(n4145), .A1N(n363), .Y(n531) );
  OAI211X2 U2377 ( .A0(n3311), .A1(n3316), .B0(n364), .C0(n531), .Y(n429) );
  CLKINVX1 U2378 ( .A(n3315), .Y(n3343) );
  BUFX20 U2379 ( .A(n4138), .Y(n3716) );
  MXI4XL U2380 ( .A(n722), .B(n877), .C(n1032), .D(n1187), .S0(n3685), .S1(
        n3715), .Y(n3345) );
  MXI4XL U2381 ( .A(n1342), .B(n1497), .C(n1652), .D(n1807), .S0(n3685), .S1(
        n3715), .Y(n3346) );
  CLKBUFX2 U2382 ( .A(n3690), .Y(n3715) );
  CLKBUFX3 U2383 ( .A(n4136), .Y(n3727) );
  MXI4XL U2384 ( .A(\CACHE[4][148] ), .B(\CACHE[5][148] ), .C(\CACHE[6][148] ), 
        .D(\CACHE[7][148] ), .S0(n3684), .S1(n3714), .Y(n3652) );
  MXI4XL U2385 ( .A(n716), .B(n871), .C(n1026), .D(n1181), .S0(n3684), .S1(
        n3714), .Y(n3347) );
  MXI4XL U2386 ( .A(n1336), .B(n1491), .C(n1646), .D(n1801), .S0(n3684), .S1(
        n3714), .Y(n3348) );
  CLKBUFX3 U2387 ( .A(n4136), .Y(n3728) );
  CLKINVX1 U2388 ( .A(n4141), .Y(n4140) );
  NAND4X2 U2389 ( .A(n547), .B(n548), .C(n549), .D(n550), .Y(n543) );
  CLKBUFX2 U2390 ( .A(n3660), .Y(n3661) );
  BUFX8 U2391 ( .A(n3659), .Y(n3663) );
  NOR2X1 U2392 ( .A(n176), .B(n7), .Y(n364) );
  NOR2X1 U2393 ( .A(n536), .B(n4141), .Y(mem_addr[0]) );
  CLKBUFX2 U2394 ( .A(n12), .Y(n4132) );
  CLKBUFX2 U2395 ( .A(n10), .Y(n4134) );
  NAND3X4 U2396 ( .A(n569), .B(n570), .C(n571), .Y(n565) );
  NAND3X4 U2397 ( .A(n562), .B(n563), .C(n564), .Y(n558) );
  NAND3X4 U2398 ( .A(n555), .B(n556), .C(n557), .Y(n551) );
  MX2X1 U2399 ( .A(n3383), .B(n3384), .S0(n3728), .Y(N34) );
  MXI4XL U2400 ( .A(n712), .B(n867), .C(n1022), .D(n1177), .S0(n3683), .S1(
        n3713), .Y(n3349) );
  MXI4XL U2401 ( .A(n1332), .B(n1487), .C(n1642), .D(n1797), .S0(n3683), .S1(
        n3713), .Y(n3350) );
  NOR2X1 U2402 ( .A(n363), .B(n533), .Y(n3351) );
  CLKBUFX2 U2403 ( .A(n3659), .Y(n3664) );
  CLKBUFX2 U2404 ( .A(n3716), .Y(n3717) );
  CLKBUFX2 U2405 ( .A(n3728), .Y(n3719) );
  CLKBUFX2 U2406 ( .A(n366), .Y(n3887) );
  NOR4X4 U2407 ( .A(n565), .B(n566), .C(n567), .D(n568), .Y(n539) );
  NOR4X4 U2408 ( .A(n558), .B(n559), .C(n560), .D(n561), .Y(n540) );
  NOR4X4 U2409 ( .A(n551), .B(n552), .C(n553), .D(n554), .Y(n541) );
  CLKBUFX2 U2410 ( .A(n433), .Y(n3881) );
  CLKBUFX2 U2411 ( .A(n467), .Y(n3876) );
  CLKBUFX2 U2412 ( .A(n353), .Y(n3892) );
  NAND3XL U2413 ( .A(n4146), .B(n3343), .C(n3351), .Y(n17) );
  NAND3BXL U2414 ( .AN(n7), .B(n8), .C(n4144), .Y(proc_stall) );
  NOR3XL U2415 ( .A(n4138), .B(n4136), .C(n4141), .Y(n349) );
  NOR3XL U2416 ( .A(n4139), .B(n4136), .C(n4141), .Y(n208) );
  NOR3XL U2417 ( .A(n4141), .B(n4138), .C(n4137), .Y(n341) );
  NOR3XL U2418 ( .A(n4141), .B(n4139), .C(n4137), .Y(n345) );
  MXI4XL U2419 ( .A(\CACHE[0][143] ), .B(\CACHE[1][143] ), .C(\CACHE[2][143] ), 
        .D(\CACHE[3][143] ), .S0(n3684), .S1(n3714), .Y(n3649) );
  MXI4XL U2420 ( .A(\CACHE[4][143] ), .B(\CACHE[5][143] ), .C(\CACHE[6][143] ), 
        .D(\CACHE[7][143] ), .S0(n3684), .S1(n3714), .Y(n3650) );
  MXI4XL U2421 ( .A(\CACHE[0][137] ), .B(\CACHE[1][137] ), .C(\CACHE[2][137] ), 
        .D(\CACHE[3][137] ), .S0(n3683), .S1(n3713), .Y(n3639) );
  MXI4XL U2422 ( .A(\CACHE[4][137] ), .B(\CACHE[5][137] ), .C(\CACHE[6][137] ), 
        .D(\CACHE[7][137] ), .S0(n3683), .S1(n3713), .Y(n3640) );
  MXI4XL U2423 ( .A(\CACHE[0][132] ), .B(\CACHE[1][132] ), .C(\CACHE[2][132] ), 
        .D(\CACHE[3][132] ), .S0(n3682), .S1(n3712), .Y(n3629) );
  MXI4XL U2424 ( .A(\CACHE[4][132] ), .B(\CACHE[5][132] ), .C(\CACHE[6][132] ), 
        .D(\CACHE[7][132] ), .S0(n3682), .S1(n3712), .Y(n3630) );
  MXI4XL U2425 ( .A(\CACHE[0][139] ), .B(\CACHE[1][139] ), .C(\CACHE[2][139] ), 
        .D(\CACHE[3][139] ), .S0(n3683), .S1(n3713), .Y(n3643) );
  MXI4XL U2426 ( .A(\CACHE[4][139] ), .B(\CACHE[5][139] ), .C(\CACHE[6][139] ), 
        .D(\CACHE[7][139] ), .S0(n3683), .S1(n3713), .Y(n3644) );
  MXI4XL U2427 ( .A(\CACHE[0][136] ), .B(\CACHE[1][136] ), .C(\CACHE[2][136] ), 
        .D(\CACHE[3][136] ), .S0(n3683), .S1(n3712), .Y(n3637) );
  MXI4XL U2428 ( .A(\CACHE[4][136] ), .B(\CACHE[5][136] ), .C(\CACHE[6][136] ), 
        .D(\CACHE[7][136] ), .S0(n3683), .S1(n3712), .Y(n3638) );
  MXI4XL U2429 ( .A(\CACHE[0][142] ), .B(\CACHE[1][142] ), .C(\CACHE[2][142] ), 
        .D(\CACHE[3][142] ), .S0(n3684), .S1(n3713), .Y(n3647) );
  MXI4XL U2430 ( .A(\CACHE[4][142] ), .B(\CACHE[5][142] ), .C(\CACHE[6][142] ), 
        .D(\CACHE[7][142] ), .S0(n3684), .S1(n3714), .Y(n3648) );
  MXI4XL U2431 ( .A(\CACHE[0][138] ), .B(\CACHE[1][138] ), .C(\CACHE[2][138] ), 
        .D(\CACHE[3][138] ), .S0(n3683), .S1(n3713), .Y(n3641) );
  MXI4XL U2432 ( .A(\CACHE[4][138] ), .B(\CACHE[5][138] ), .C(\CACHE[6][138] ), 
        .D(\CACHE[7][138] ), .S0(n3683), .S1(n3714), .Y(n3642) );
  MXI4XL U2433 ( .A(\CACHE[0][141] ), .B(\CACHE[1][141] ), .C(\CACHE[2][141] ), 
        .D(\CACHE[3][141] ), .S0(n3683), .S1(n3713), .Y(n3645) );
  MXI4XL U2434 ( .A(\CACHE[4][141] ), .B(\CACHE[5][141] ), .C(\CACHE[6][141] ), 
        .D(\CACHE[7][141] ), .S0(n3683), .S1(n3713), .Y(n3646) );
  MX4XL U2435 ( .A(\CACHE[0][128] ), .B(\CACHE[1][128] ), .C(\CACHE[2][128] ), 
        .D(\CACHE[3][128] ), .S0(n3681), .S1(n3711), .Y(n3352) );
  MX4XL U2436 ( .A(\CACHE[4][128] ), .B(\CACHE[5][128] ), .C(\CACHE[6][128] ), 
        .D(\CACHE[7][128] ), .S0(n3660), .S1(n3711), .Y(n3353) );
  MX4XL U2437 ( .A(n724), .B(n879), .C(n1034), .D(n1189), .S0(n3685), .S1(
        n3718), .Y(n3655) );
  MX4XL U2438 ( .A(n1344), .B(n1499), .C(n1654), .D(n1809), .S0(n3685), .S1(
        n3716), .Y(n3656) );
  MX4XL U2439 ( .A(n705), .B(n860), .C(n1015), .D(n1170), .S0(n3682), .S1(
        n3712), .Y(n3631) );
  MX4XL U2440 ( .A(n1325), .B(n1480), .C(n1635), .D(n1790), .S0(n3682), .S1(
        n3712), .Y(n3632) );
  MX4XL U2441 ( .A(n1327), .B(n1482), .C(n1637), .D(n1792), .S0(n3682), .S1(
        n3712), .Y(n3636) );
  MX4XL U2442 ( .A(n706), .B(n861), .C(n1016), .D(n1171), .S0(n3682), .S1(
        n3712), .Y(n3633) );
  MX4XL U2443 ( .A(n1326), .B(n1481), .C(n1636), .D(n1791), .S0(n3682), .S1(
        n3712), .Y(n3634) );
  XNOR2X4 U2444 ( .A(N51), .B(proc_addr[13]), .Y(n555) );
  XNOR2X4 U2445 ( .A(N55), .B(proc_addr[9]), .Y(n556) );
  XNOR2X4 U2446 ( .A(N46), .B(proc_addr[18]), .Y(n557) );
  XNOR2X4 U2447 ( .A(N48), .B(proc_addr[16]), .Y(n569) );
  XNOR2X4 U2448 ( .A(N49), .B(proc_addr[15]), .Y(n570) );
  XNOR2X4 U2449 ( .A(N38), .B(proc_addr[26]), .Y(n571) );
  MX4XL U2450 ( .A(n702), .B(n857), .C(n1012), .D(n1167), .S0(n3682), .S1(
        n3711), .Y(n3625) );
  MX4XL U2451 ( .A(n1322), .B(n1477), .C(n1632), .D(n1787), .S0(n3682), .S1(
        n3711), .Y(n3626) );
  NAND2BXL U2452 ( .AN(N33), .B(n3317), .Y(n8) );
  NAND3XL U2453 ( .A(n3351), .B(n4146), .C(n3315), .Y(n12) );
  NAND3XL U2454 ( .A(n3351), .B(n3343), .C(n3313), .Y(n10) );
  NAND3XL U2455 ( .A(n3313), .B(n3351), .C(n3315), .Y(n15) );
  MX4XL U2456 ( .A(\CACHE[0][153] ), .B(\CACHE[1][153] ), .C(\CACHE[2][153] ), 
        .D(\CACHE[3][153] ), .S0(n3685), .S1(n3715), .Y(n3383) );
  MX4XL U2457 ( .A(\CACHE[4][153] ), .B(\CACHE[5][153] ), .C(\CACHE[6][153] ), 
        .D(\CACHE[7][153] ), .S0(n3685), .S1(n3715), .Y(n3384) );
  MX4XL U2458 ( .A(n726), .B(n881), .C(n1036), .D(n1191), .S0(n3685), .S1(
        n3715), .Y(n3657) );
  MX4XL U2459 ( .A(n1346), .B(n1501), .C(n1656), .D(n1811), .S0(n3685), .S1(
        n3715), .Y(n3658) );
  AND2XL U2460 ( .A(n364), .B(n3311), .Y(n362) );
  NAND4BXL U2461 ( .AN(n3311), .B(N34), .C(n537), .D(n533), .Y(n535) );
  OAI2BB1XL U2462 ( .A0N(n3316), .A1N(proc_write), .B0(n363), .Y(n537) );
  OAI211XL U2463 ( .A0(n359), .A1(n4145), .B0(n361), .C0(n362), .Y(n358) );
  AND2XL U2464 ( .A(n363), .B(n3317), .Y(n359) );
  NOR2X1 U2465 ( .A(n3317), .B(proc_write), .Y(n7) );
  MXI2X1 U2466 ( .A(n3355), .B(n3356), .S0(n3726), .Y(n3354) );
  MX4X1 U2467 ( .A(\CACHE[0][119] ), .B(\CACHE[1][119] ), .C(\CACHE[2][119] ), 
        .D(\CACHE[3][119] ), .S0(n3680), .S1(n3694), .Y(n3355) );
  MX4X1 U2468 ( .A(\CACHE[4][119] ), .B(\CACHE[5][119] ), .C(\CACHE[6][119] ), 
        .D(\CACHE[7][119] ), .S0(n3680), .S1(n3696), .Y(n3356) );
  MXI2X1 U2469 ( .A(n3358), .B(n3359), .S0(n3726), .Y(n3357) );
  MX4X1 U2470 ( .A(\CACHE[0][120] ), .B(\CACHE[1][120] ), .C(\CACHE[2][120] ), 
        .D(\CACHE[3][120] ), .S0(n3680), .S1(n3693), .Y(n3358) );
  MX4X1 U2471 ( .A(\CACHE[4][120] ), .B(\CACHE[5][120] ), .C(\CACHE[6][120] ), 
        .D(\CACHE[7][120] ), .S0(n3680), .S1(n3697), .Y(n3359) );
  MXI2X1 U2472 ( .A(n3361), .B(n3362), .S0(n3726), .Y(n3360) );
  MX4X1 U2473 ( .A(\CACHE[0][121] ), .B(\CACHE[1][121] ), .C(\CACHE[2][121] ), 
        .D(\CACHE[3][121] ), .S0(n3680), .S1(n3687), .Y(n3361) );
  MX4X1 U2474 ( .A(\CACHE[4][121] ), .B(\CACHE[5][121] ), .C(\CACHE[6][121] ), 
        .D(\CACHE[7][121] ), .S0(n3680), .S1(n3706), .Y(n3362) );
  MXI2X1 U2475 ( .A(n3364), .B(n3365), .S0(n3726), .Y(n3363) );
  MX4XL U2476 ( .A(\CACHE[0][122] ), .B(\CACHE[1][122] ), .C(\CACHE[2][122] ), 
        .D(\CACHE[3][122] ), .S0(n3681), .S1(n3696), .Y(n3364) );
  MX4X1 U2477 ( .A(\CACHE[4][122] ), .B(\CACHE[5][122] ), .C(\CACHE[6][122] ), 
        .D(\CACHE[7][122] ), .S0(n3680), .S1(n3687), .Y(n3365) );
  MXI2X1 U2478 ( .A(n3367), .B(n3368), .S0(n3726), .Y(n3366) );
  MX4XL U2479 ( .A(\CACHE[0][123] ), .B(\CACHE[1][123] ), .C(\CACHE[2][123] ), 
        .D(\CACHE[3][123] ), .S0(n3681), .S1(n3696), .Y(n3367) );
  MX4XL U2480 ( .A(\CACHE[4][123] ), .B(\CACHE[5][123] ), .C(\CACHE[6][123] ), 
        .D(\CACHE[7][123] ), .S0(n3681), .S1(n3694), .Y(n3368) );
  MXI2X1 U2481 ( .A(n3370), .B(n3371), .S0(n3726), .Y(n3369) );
  MX4XL U2482 ( .A(\CACHE[0][124] ), .B(\CACHE[1][124] ), .C(\CACHE[2][124] ), 
        .D(\CACHE[3][124] ), .S0(n3681), .S1(n3709), .Y(n3370) );
  MX4XL U2483 ( .A(\CACHE[4][124] ), .B(\CACHE[5][124] ), .C(\CACHE[6][124] ), 
        .D(\CACHE[7][124] ), .S0(n3681), .S1(n3708), .Y(n3371) );
  MXI2X1 U2484 ( .A(n3373), .B(n3374), .S0(n3726), .Y(n3372) );
  MX4XL U2485 ( .A(\CACHE[0][125] ), .B(\CACHE[1][125] ), .C(\CACHE[2][125] ), 
        .D(\CACHE[3][125] ), .S0(n3681), .S1(n3711), .Y(n3373) );
  MX4XL U2486 ( .A(\CACHE[4][125] ), .B(\CACHE[5][125] ), .C(\CACHE[6][125] ), 
        .D(\CACHE[7][125] ), .S0(n3681), .S1(n3711), .Y(n3374) );
  MXI2X1 U2487 ( .A(n3376), .B(n3377), .S0(n3726), .Y(n3375) );
  MX4XL U2488 ( .A(\CACHE[0][126] ), .B(\CACHE[1][126] ), .C(\CACHE[2][126] ), 
        .D(\CACHE[3][126] ), .S0(n3681), .S1(n3711), .Y(n3376) );
  MX4XL U2489 ( .A(\CACHE[4][126] ), .B(\CACHE[5][126] ), .C(\CACHE[6][126] ), 
        .D(\CACHE[7][126] ), .S0(n3681), .S1(n3711), .Y(n3377) );
  MXI2X1 U2490 ( .A(n3379), .B(n3380), .S0(n3726), .Y(n3378) );
  MX4XL U2491 ( .A(\CACHE[0][127] ), .B(\CACHE[1][127] ), .C(\CACHE[2][127] ), 
        .D(\CACHE[3][127] ), .S0(n3681), .S1(n3711), .Y(n3379) );
  MX4XL U2492 ( .A(\CACHE[4][127] ), .B(\CACHE[5][127] ), .C(\CACHE[6][127] ), 
        .D(\CACHE[7][127] ), .S0(n3681), .S1(n3711), .Y(n3380) );
  CLKINVX1 U2493 ( .A(proc_wdata[0]), .Y(n4178) );
  CLKINVX1 U2494 ( .A(proc_wdata[1]), .Y(n4177) );
  CLKINVX1 U2495 ( .A(proc_wdata[2]), .Y(n4176) );
  CLKINVX1 U2496 ( .A(proc_wdata[3]), .Y(n4175) );
  CLKINVX1 U2497 ( .A(proc_wdata[4]), .Y(n4174) );
  CLKINVX1 U2498 ( .A(proc_wdata[5]), .Y(n4173) );
  CLKINVX1 U2499 ( .A(proc_wdata[6]), .Y(n4172) );
  CLKINVX1 U2500 ( .A(proc_wdata[7]), .Y(n4171) );
  CLKINVX1 U2501 ( .A(proc_wdata[8]), .Y(n4170) );
  CLKINVX1 U2502 ( .A(proc_wdata[9]), .Y(n4169) );
  CLKINVX1 U2503 ( .A(proc_wdata[10]), .Y(n4168) );
  CLKINVX1 U2504 ( .A(proc_wdata[11]), .Y(n4167) );
  CLKINVX1 U2505 ( .A(proc_wdata[12]), .Y(n4166) );
  CLKINVX1 U2506 ( .A(proc_wdata[13]), .Y(n4165) );
  CLKINVX1 U2507 ( .A(proc_wdata[14]), .Y(n4164) );
  CLKINVX1 U2508 ( .A(proc_wdata[15]), .Y(n4163) );
  CLKINVX1 U2509 ( .A(proc_wdata[16]), .Y(n4162) );
  CLKINVX1 U2510 ( .A(proc_wdata[17]), .Y(n4161) );
  CLKINVX1 U2511 ( .A(proc_wdata[18]), .Y(n4160) );
  CLKINVX1 U2512 ( .A(proc_wdata[19]), .Y(n4159) );
  CLKINVX1 U2513 ( .A(proc_wdata[20]), .Y(n4158) );
  CLKINVX1 U2514 ( .A(proc_wdata[21]), .Y(n4157) );
  CLKINVX1 U2515 ( .A(proc_wdata[22]), .Y(n4156) );
  CLKINVX1 U2516 ( .A(proc_wdata[23]), .Y(n4155) );
  CLKINVX1 U2517 ( .A(proc_wdata[24]), .Y(n4154) );
  CLKINVX1 U2518 ( .A(proc_wdata[25]), .Y(n4153) );
  CLKINVX1 U2519 ( .A(proc_wdata[26]), .Y(n4152) );
  CLKINVX1 U2520 ( .A(proc_wdata[27]), .Y(n4151) );
  CLKINVX1 U2521 ( .A(proc_wdata[28]), .Y(n4150) );
  CLKINVX1 U2522 ( .A(proc_wdata[29]), .Y(n4149) );
  CLKINVX1 U2523 ( .A(proc_wdata[30]), .Y(n4148) );
  CLKINVX1 U2524 ( .A(proc_wdata[31]), .Y(n4147) );
  AOI22X2 U2525 ( .A0(n3889), .A1(n3245), .B0(proc_addr[25]), .B1(n3901), .Y(
        n201) );
  XNOR2X1 U2526 ( .A(n3245), .B(proc_addr[25]), .Y(n547) );
  MXI4XL U2527 ( .A(\CACHE[0][148] ), .B(\CACHE[1][148] ), .C(\CACHE[2][148] ), 
        .D(\CACHE[3][148] ), .S0(n3685), .S1(n3714), .Y(n3651) );
  CLKBUFX3 U2528 ( .A(n3692), .Y(n3711) );
  INVX3 U2529 ( .A(n3944), .Y(n3932) );
  INVX3 U2530 ( .A(n3944), .Y(n3933) );
  INVX3 U2531 ( .A(n3947), .Y(n3934) );
  INVX3 U2532 ( .A(n3944), .Y(n3935) );
  INVX3 U2533 ( .A(n3955), .Y(n3936) );
  INVX3 U2534 ( .A(n3944), .Y(n3937) );
  INVX3 U2535 ( .A(n3944), .Y(n3938) );
  INVX3 U2536 ( .A(n3944), .Y(n3939) );
  INVX3 U2537 ( .A(n3944), .Y(n3940) );
  INVX3 U2538 ( .A(n3946), .Y(n3941) );
  INVX3 U2539 ( .A(n3945), .Y(n3942) );
  INVX3 U2540 ( .A(n3945), .Y(n3931) );
  INVX3 U2541 ( .A(n3952), .Y(n3943) );
  CLKBUFX3 U2542 ( .A(n3694), .Y(n3698) );
  CLKBUFX3 U2543 ( .A(n3686), .Y(n3699) );
  CLKBUFX3 U2544 ( .A(n3686), .Y(n3700) );
  CLKBUFX3 U2545 ( .A(n3695), .Y(n3701) );
  CLKBUFX3 U2546 ( .A(n3694), .Y(n3702) );
  CLKBUFX3 U2547 ( .A(n3695), .Y(n3703) );
  CLKBUFX3 U2548 ( .A(n3695), .Y(n3704) );
  CLKBUFX3 U2549 ( .A(n3695), .Y(n3705) );
  CLKBUFX3 U2550 ( .A(n3694), .Y(n3706) );
  CLKBUFX3 U2551 ( .A(n3694), .Y(n3707) );
  CLKBUFX3 U2552 ( .A(n3693), .Y(n3708) );
  CLKBUFX3 U2553 ( .A(n3693), .Y(n3709) );
  CLKBUFX3 U2554 ( .A(n3687), .Y(n3710) );
  CLKBUFX3 U2555 ( .A(n4136), .Y(n3726) );
  CLKBUFX3 U2556 ( .A(n3662), .Y(n3682) );
  CLKBUFX3 U2557 ( .A(n3662), .Y(n3683) );
  CLKBUFX3 U2558 ( .A(n3661), .Y(n3684) );
  CLKBUFX3 U2559 ( .A(n3661), .Y(n3685) );
  CLKBUFX3 U2560 ( .A(n3689), .Y(n3691) );
  CLKBUFX3 U2561 ( .A(n3689), .Y(n3690) );
  CLKBUFX3 U2562 ( .A(n3719), .Y(n3721) );
  CLKBUFX3 U2563 ( .A(n3719), .Y(n3722) );
  CLKBUFX3 U2564 ( .A(n3719), .Y(n3723) );
  CLKBUFX3 U2565 ( .A(n3719), .Y(n3724) );
  CLKBUFX3 U2566 ( .A(n3719), .Y(n3725) );
  CLKBUFX3 U2567 ( .A(n3664), .Y(n3666) );
  CLKBUFX3 U2568 ( .A(n3664), .Y(n3667) );
  CLKBUFX3 U2569 ( .A(n3665), .Y(n3668) );
  CLKBUFX3 U2570 ( .A(n3664), .Y(n3669) );
  CLKBUFX3 U2571 ( .A(n3664), .Y(n3670) );
  CLKBUFX3 U2572 ( .A(n3665), .Y(n3671) );
  CLKBUFX3 U2573 ( .A(n3664), .Y(n3672) );
  CLKBUFX3 U2574 ( .A(n3665), .Y(n3673) );
  CLKBUFX3 U2575 ( .A(n3664), .Y(n3674) );
  CLKBUFX3 U2576 ( .A(n3664), .Y(n3675) );
  CLKBUFX3 U2577 ( .A(n3664), .Y(n3676) );
  CLKBUFX3 U2578 ( .A(n3664), .Y(n3677) );
  CLKBUFX3 U2579 ( .A(n3664), .Y(n3678) );
  CLKBUFX3 U2580 ( .A(n3664), .Y(n3679) );
  CLKBUFX3 U2581 ( .A(n3663), .Y(n3680) );
  CLKBUFX3 U2582 ( .A(n3957), .Y(n3944) );
  CLKBUFX3 U2583 ( .A(n3957), .Y(n3945) );
  CLKBUFX3 U2584 ( .A(n3957), .Y(n3946) );
  CLKBUFX3 U2585 ( .A(n3958), .Y(n3948) );
  CLKBUFX3 U2586 ( .A(n3958), .Y(n3949) );
  CLKBUFX3 U2587 ( .A(n3958), .Y(n3950) );
  CLKBUFX3 U2588 ( .A(n3958), .Y(n3951) );
  CLKBUFX3 U2589 ( .A(n3957), .Y(n3952) );
  CLKBUFX3 U2590 ( .A(n3957), .Y(n3953) );
  CLKBUFX3 U2591 ( .A(n3945), .Y(n3954) );
  CLKBUFX3 U2592 ( .A(n3957), .Y(n3955) );
  CLKBUFX3 U2593 ( .A(n3944), .Y(n3956) );
  INVX3 U2594 ( .A(n3926), .Y(n3904) );
  INVX3 U2595 ( .A(n3927), .Y(n3905) );
  INVX3 U2596 ( .A(n3928), .Y(n3906) );
  INVX3 U2597 ( .A(n3916), .Y(n3907) );
  INVX3 U2598 ( .A(n3916), .Y(n3908) );
  INVX3 U2599 ( .A(n3917), .Y(n3909) );
  INVX3 U2600 ( .A(n3929), .Y(n3910) );
  INVX3 U2601 ( .A(n3929), .Y(n3911) );
  INVX3 U2602 ( .A(n3928), .Y(n3912) );
  INVX3 U2603 ( .A(n3927), .Y(n3913) );
  INVX3 U2604 ( .A(n3917), .Y(n3914) );
  INVX3 U2605 ( .A(n4114), .Y(n4102) );
  INVX3 U2606 ( .A(n4111), .Y(n4103) );
  INVX3 U2607 ( .A(n4116), .Y(n4104) );
  INVX3 U2608 ( .A(n4112), .Y(n4105) );
  INVX3 U2609 ( .A(n4111), .Y(n4106) );
  INVX3 U2610 ( .A(n4112), .Y(n4107) );
  INVX3 U2611 ( .A(n4111), .Y(n4108) );
  INVX3 U2612 ( .A(n4111), .Y(n4109) );
  INVX3 U2613 ( .A(n4111), .Y(n4110) );
  INVX3 U2614 ( .A(n4111), .Y(n4100) );
  INVX3 U2615 ( .A(n4114), .Y(n4101) );
  INVX3 U2616 ( .A(n4094), .Y(n4072) );
  INVX3 U2617 ( .A(n4095), .Y(n4073) );
  INVX3 U2618 ( .A(n4096), .Y(n4074) );
  INVX3 U2619 ( .A(n4084), .Y(n4075) );
  INVX3 U2620 ( .A(n4084), .Y(n4076) );
  INVX3 U2621 ( .A(n4085), .Y(n4077) );
  INVX3 U2622 ( .A(n4097), .Y(n4078) );
  INVX3 U2623 ( .A(n4097), .Y(n4079) );
  INVX3 U2624 ( .A(n4096), .Y(n4080) );
  INVX3 U2625 ( .A(n4095), .Y(n4081) );
  INVX3 U2626 ( .A(n4085), .Y(n4082) );
  INVX3 U2627 ( .A(n4066), .Y(n4044) );
  INVX3 U2628 ( .A(n4055), .Y(n4045) );
  INVX3 U2629 ( .A(n4062), .Y(n4046) );
  INVX3 U2630 ( .A(n4056), .Y(n4047) );
  INVX3 U2631 ( .A(n4064), .Y(n4048) );
  INVX3 U2632 ( .A(n4055), .Y(n4049) );
  INVX3 U2633 ( .A(n4055), .Y(n4050) );
  INVX3 U2634 ( .A(n4055), .Y(n4051) );
  INVX3 U2635 ( .A(n4055), .Y(n4052) );
  INVX3 U2636 ( .A(n4055), .Y(n4053) );
  INVX3 U2637 ( .A(n4055), .Y(n4054) );
  INVX3 U2638 ( .A(n4038), .Y(n4016) );
  INVX3 U2639 ( .A(n4039), .Y(n4017) );
  INVX3 U2640 ( .A(n4040), .Y(n4018) );
  INVX3 U2641 ( .A(n4028), .Y(n4019) );
  INVX3 U2642 ( .A(n4028), .Y(n4020) );
  INVX3 U2643 ( .A(n4029), .Y(n4021) );
  INVX3 U2644 ( .A(n4041), .Y(n4022) );
  INVX3 U2645 ( .A(n4041), .Y(n4023) );
  INVX3 U2646 ( .A(n4040), .Y(n4024) );
  INVX3 U2647 ( .A(n4039), .Y(n4025) );
  INVX3 U2648 ( .A(n4029), .Y(n4026) );
  INVX3 U2649 ( .A(n4010), .Y(n3988) );
  INVX3 U2650 ( .A(n3999), .Y(n3989) );
  INVX3 U2651 ( .A(n4006), .Y(n3990) );
  INVX3 U2652 ( .A(n4000), .Y(n3991) );
  INVX3 U2653 ( .A(n4008), .Y(n3992) );
  INVX3 U2654 ( .A(n3999), .Y(n3993) );
  INVX3 U2655 ( .A(n3999), .Y(n3994) );
  INVX3 U2656 ( .A(n3999), .Y(n3995) );
  INVX3 U2657 ( .A(n3999), .Y(n3996) );
  INVX3 U2658 ( .A(n3999), .Y(n3997) );
  INVX3 U2659 ( .A(n3999), .Y(n3998) );
  INVX3 U2660 ( .A(n3982), .Y(n3960) );
  INVX3 U2661 ( .A(n3983), .Y(n3961) );
  INVX3 U2662 ( .A(n3984), .Y(n3962) );
  INVX3 U2663 ( .A(n3972), .Y(n3963) );
  INVX3 U2664 ( .A(n3972), .Y(n3964) );
  INVX3 U2665 ( .A(n3973), .Y(n3965) );
  INVX3 U2666 ( .A(n3985), .Y(n3966) );
  INVX3 U2667 ( .A(n3985), .Y(n3967) );
  INVX3 U2668 ( .A(n3984), .Y(n3968) );
  INVX3 U2669 ( .A(n3983), .Y(n3969) );
  INVX3 U2670 ( .A(n3973), .Y(n3970) );
  INVX3 U2671 ( .A(n3916), .Y(n3903) );
  INVX3 U2672 ( .A(n4112), .Y(n4099) );
  INVX3 U2673 ( .A(n4084), .Y(n4071) );
  INVX3 U2674 ( .A(n4058), .Y(n4043) );
  INVX3 U2675 ( .A(n4028), .Y(n4015) );
  INVX3 U2676 ( .A(n4002), .Y(n3987) );
  INVX3 U2677 ( .A(n3972), .Y(n3959) );
  CLKBUFX3 U2678 ( .A(n3664), .Y(n3665) );
  INVX3 U2679 ( .A(n3926), .Y(n3915) );
  INVX3 U2680 ( .A(n4094), .Y(n4083) );
  INVX3 U2681 ( .A(n4038), .Y(n4027) );
  INVX3 U2682 ( .A(n3982), .Y(n3971) );
  CLKBUFX3 U2683 ( .A(n3717), .Y(n3695) );
  CLKBUFX3 U2684 ( .A(n3717), .Y(n3694) );
  CLKBUFX3 U2685 ( .A(n3687), .Y(n3693) );
  CLKBUFX3 U2686 ( .A(n3718), .Y(n3688) );
  CLKBUFX3 U2687 ( .A(n3660), .Y(n3662) );
  CLKBUFX3 U2688 ( .A(n3719), .Y(n3720) );
  CLKBUFX3 U2689 ( .A(n4121), .Y(n4111) );
  CLKBUFX3 U2690 ( .A(n4057), .Y(n4055) );
  CLKBUFX3 U2691 ( .A(n4001), .Y(n3999) );
  CLKBUFX3 U2692 ( .A(n3930), .Y(n3916) );
  CLKBUFX3 U2693 ( .A(n4120), .Y(n4112) );
  CLKBUFX3 U2694 ( .A(n4098), .Y(n4084) );
  CLKBUFX3 U2695 ( .A(n4042), .Y(n4028) );
  CLKBUFX3 U2696 ( .A(n3986), .Y(n3972) );
  CLKBUFX3 U2697 ( .A(n3930), .Y(n3917) );
  CLKBUFX3 U2698 ( .A(n3929), .Y(n3918) );
  CLKBUFX3 U2699 ( .A(n3916), .Y(n3919) );
  CLKBUFX3 U2700 ( .A(n3929), .Y(n3920) );
  CLKBUFX3 U2701 ( .A(n3929), .Y(n3921) );
  CLKBUFX3 U2702 ( .A(n3929), .Y(n3922) );
  CLKBUFX3 U2703 ( .A(n3929), .Y(n3923) );
  CLKBUFX3 U2704 ( .A(n3929), .Y(n3924) );
  CLKBUFX3 U2705 ( .A(n3919), .Y(n3925) );
  CLKBUFX3 U2706 ( .A(n3930), .Y(n3926) );
  CLKBUFX3 U2707 ( .A(n3930), .Y(n3927) );
  CLKBUFX3 U2708 ( .A(n3930), .Y(n3928) );
  CLKBUFX3 U2709 ( .A(n4125), .Y(n4115) );
  CLKBUFX3 U2710 ( .A(n4125), .Y(n4116) );
  CLKBUFX3 U2711 ( .A(n4125), .Y(n4117) );
  CLKBUFX3 U2712 ( .A(n4125), .Y(n4118) );
  CLKBUFX3 U2713 ( .A(n4125), .Y(n4119) );
  CLKBUFX3 U2714 ( .A(n4126), .Y(n4120) );
  CLKBUFX3 U2715 ( .A(n4126), .Y(n4121) );
  CLKBUFX3 U2716 ( .A(n4126), .Y(n4122) );
  CLKBUFX3 U2717 ( .A(n4126), .Y(n4123) );
  CLKBUFX3 U2718 ( .A(n4126), .Y(n4124) );
  CLKBUFX3 U2719 ( .A(n4122), .Y(n4113) );
  CLKBUFX3 U2720 ( .A(n4098), .Y(n4085) );
  CLKBUFX3 U2721 ( .A(n4097), .Y(n4086) );
  CLKBUFX3 U2722 ( .A(n4084), .Y(n4087) );
  CLKBUFX3 U2723 ( .A(n4097), .Y(n4088) );
  CLKBUFX3 U2724 ( .A(n4097), .Y(n4089) );
  CLKBUFX3 U2725 ( .A(n4097), .Y(n4090) );
  CLKBUFX3 U2726 ( .A(n4097), .Y(n4091) );
  CLKBUFX3 U2727 ( .A(n4097), .Y(n4092) );
  CLKBUFX3 U2728 ( .A(n4087), .Y(n4093) );
  CLKBUFX3 U2729 ( .A(n4098), .Y(n4094) );
  CLKBUFX3 U2730 ( .A(n4098), .Y(n4095) );
  CLKBUFX3 U2731 ( .A(n4098), .Y(n4096) );
  CLKBUFX3 U2732 ( .A(n4061), .Y(n4056) );
  CLKBUFX3 U2733 ( .A(n4069), .Y(n4057) );
  CLKBUFX3 U2734 ( .A(n4069), .Y(n4058) );
  CLKBUFX3 U2735 ( .A(n4069), .Y(n4059) );
  CLKBUFX3 U2736 ( .A(n4069), .Y(n4060) );
  CLKBUFX3 U2737 ( .A(n4069), .Y(n4061) );
  CLKBUFX3 U2738 ( .A(n4069), .Y(n4062) );
  CLKBUFX3 U2739 ( .A(n4070), .Y(n4063) );
  CLKBUFX3 U2740 ( .A(n4070), .Y(n4064) );
  CLKBUFX3 U2741 ( .A(n4070), .Y(n4065) );
  CLKBUFX3 U2742 ( .A(n4070), .Y(n4066) );
  CLKBUFX3 U2743 ( .A(n4070), .Y(n4067) );
  CLKBUFX3 U2744 ( .A(n4070), .Y(n4068) );
  CLKBUFX3 U2745 ( .A(n4042), .Y(n4029) );
  CLKBUFX3 U2746 ( .A(n4041), .Y(n4030) );
  CLKBUFX3 U2747 ( .A(n4028), .Y(n4031) );
  CLKBUFX3 U2748 ( .A(n4041), .Y(n4032) );
  CLKBUFX3 U2749 ( .A(n4041), .Y(n4033) );
  CLKBUFX3 U2750 ( .A(n4041), .Y(n4034) );
  CLKBUFX3 U2751 ( .A(n4041), .Y(n4035) );
  CLKBUFX3 U2752 ( .A(n4041), .Y(n4036) );
  CLKBUFX3 U2753 ( .A(n4031), .Y(n4037) );
  CLKBUFX3 U2754 ( .A(n4042), .Y(n4038) );
  CLKBUFX3 U2755 ( .A(n4042), .Y(n4039) );
  CLKBUFX3 U2756 ( .A(n4042), .Y(n4040) );
  CLKBUFX3 U2757 ( .A(n4005), .Y(n4000) );
  CLKBUFX3 U2758 ( .A(n4013), .Y(n4001) );
  CLKBUFX3 U2759 ( .A(n4013), .Y(n4002) );
  CLKBUFX3 U2760 ( .A(n4013), .Y(n4003) );
  CLKBUFX3 U2761 ( .A(n4013), .Y(n4004) );
  CLKBUFX3 U2762 ( .A(n4013), .Y(n4005) );
  CLKBUFX3 U2763 ( .A(n4013), .Y(n4006) );
  CLKBUFX3 U2764 ( .A(n4014), .Y(n4007) );
  CLKBUFX3 U2765 ( .A(n4014), .Y(n4008) );
  CLKBUFX3 U2766 ( .A(n4014), .Y(n4009) );
  CLKBUFX3 U2767 ( .A(n4014), .Y(n4010) );
  CLKBUFX3 U2768 ( .A(n4014), .Y(n4011) );
  CLKBUFX3 U2769 ( .A(n4014), .Y(n4012) );
  CLKBUFX3 U2770 ( .A(n3986), .Y(n3973) );
  CLKBUFX3 U2771 ( .A(n3985), .Y(n3974) );
  CLKBUFX3 U2772 ( .A(n3972), .Y(n3975) );
  CLKBUFX3 U2773 ( .A(n3985), .Y(n3976) );
  CLKBUFX3 U2774 ( .A(n3985), .Y(n3977) );
  CLKBUFX3 U2775 ( .A(n3985), .Y(n3978) );
  CLKBUFX3 U2776 ( .A(n3985), .Y(n3979) );
  CLKBUFX3 U2777 ( .A(n3985), .Y(n3980) );
  CLKBUFX3 U2778 ( .A(n3975), .Y(n3981) );
  CLKBUFX3 U2779 ( .A(n3986), .Y(n3982) );
  CLKBUFX3 U2780 ( .A(n3986), .Y(n3983) );
  CLKBUFX3 U2781 ( .A(n3986), .Y(n3984) );
  CLKBUFX3 U2782 ( .A(n3686), .Y(n3697) );
  CLKBUFX3 U2783 ( .A(n3695), .Y(n3696) );
  CLKBUFX3 U2784 ( .A(n3717), .Y(n3686) );
  CLKBUFX3 U2785 ( .A(n3718), .Y(n3687) );
  CLKBUFX3 U2786 ( .A(n3860), .Y(n3734) );
  CLKBUFX3 U2787 ( .A(n3860), .Y(n3735) );
  CLKBUFX3 U2788 ( .A(n3860), .Y(n3736) );
  CLKBUFX3 U2789 ( .A(n3860), .Y(n3737) );
  CLKBUFX3 U2790 ( .A(n3859), .Y(n3738) );
  CLKBUFX3 U2791 ( .A(n3859), .Y(n3739) );
  CLKBUFX3 U2792 ( .A(n3859), .Y(n3740) );
  CLKBUFX3 U2793 ( .A(n3859), .Y(n3741) );
  CLKBUFX3 U2794 ( .A(n3858), .Y(n3742) );
  CLKBUFX3 U2795 ( .A(n3858), .Y(n3743) );
  CLKBUFX3 U2796 ( .A(n3858), .Y(n3744) );
  CLKBUFX3 U2797 ( .A(n3858), .Y(n3745) );
  CLKBUFX3 U2798 ( .A(n3857), .Y(n3746) );
  CLKBUFX3 U2799 ( .A(n3857), .Y(n3747) );
  CLKBUFX3 U2800 ( .A(n3857), .Y(n3748) );
  CLKBUFX3 U2801 ( .A(n3857), .Y(n3749) );
  CLKBUFX3 U2802 ( .A(n3856), .Y(n3750) );
  CLKBUFX3 U2803 ( .A(n3856), .Y(n3751) );
  CLKBUFX3 U2804 ( .A(n3856), .Y(n3752) );
  CLKBUFX3 U2805 ( .A(n3856), .Y(n3753) );
  CLKBUFX3 U2806 ( .A(n3855), .Y(n3754) );
  CLKBUFX3 U2807 ( .A(n3855), .Y(n3755) );
  CLKBUFX3 U2808 ( .A(n3855), .Y(n3756) );
  CLKBUFX3 U2809 ( .A(n3855), .Y(n3757) );
  CLKBUFX3 U2810 ( .A(n3854), .Y(n3758) );
  CLKBUFX3 U2811 ( .A(n3854), .Y(n3759) );
  CLKBUFX3 U2812 ( .A(n3854), .Y(n3760) );
  CLKBUFX3 U2813 ( .A(n3854), .Y(n3761) );
  CLKBUFX3 U2814 ( .A(n3853), .Y(n3762) );
  CLKBUFX3 U2815 ( .A(n3853), .Y(n3763) );
  CLKBUFX3 U2816 ( .A(n3853), .Y(n3764) );
  CLKBUFX3 U2817 ( .A(n3853), .Y(n3765) );
  CLKBUFX3 U2818 ( .A(n3852), .Y(n3766) );
  CLKBUFX3 U2819 ( .A(n3852), .Y(n3767) );
  CLKBUFX3 U2820 ( .A(n3852), .Y(n3768) );
  CLKBUFX3 U2821 ( .A(n3852), .Y(n3769) );
  CLKBUFX3 U2822 ( .A(n3851), .Y(n3770) );
  CLKBUFX3 U2823 ( .A(n3851), .Y(n3771) );
  CLKBUFX3 U2824 ( .A(n3851), .Y(n3772) );
  CLKBUFX3 U2825 ( .A(n3851), .Y(n3773) );
  CLKBUFX3 U2826 ( .A(n3850), .Y(n3774) );
  CLKBUFX3 U2827 ( .A(n3850), .Y(n3775) );
  CLKBUFX3 U2828 ( .A(n3850), .Y(n3776) );
  CLKBUFX3 U2829 ( .A(n3850), .Y(n3777) );
  CLKBUFX3 U2830 ( .A(n3849), .Y(n3778) );
  CLKBUFX3 U2831 ( .A(n3849), .Y(n3779) );
  CLKBUFX3 U2832 ( .A(n3849), .Y(n3780) );
  CLKBUFX3 U2833 ( .A(n3849), .Y(n3781) );
  CLKBUFX3 U2834 ( .A(n3732), .Y(n3782) );
  CLKBUFX3 U2835 ( .A(n3732), .Y(n3783) );
  CLKBUFX3 U2836 ( .A(n3842), .Y(n3784) );
  CLKBUFX3 U2837 ( .A(n3838), .Y(n3785) );
  CLKBUFX3 U2838 ( .A(n3848), .Y(n3786) );
  CLKBUFX3 U2839 ( .A(n3848), .Y(n3787) );
  CLKBUFX3 U2840 ( .A(n3848), .Y(n3788) );
  CLKBUFX3 U2841 ( .A(n3848), .Y(n3789) );
  CLKBUFX3 U2842 ( .A(n3847), .Y(n3790) );
  CLKBUFX3 U2843 ( .A(n3847), .Y(n3791) );
  CLKBUFX3 U2844 ( .A(n3847), .Y(n3792) );
  CLKBUFX3 U2845 ( .A(n3847), .Y(n3793) );
  CLKBUFX3 U2846 ( .A(n3846), .Y(n3794) );
  CLKBUFX3 U2847 ( .A(n3846), .Y(n3795) );
  CLKBUFX3 U2848 ( .A(n3846), .Y(n3796) );
  CLKBUFX3 U2849 ( .A(n3846), .Y(n3797) );
  CLKBUFX3 U2850 ( .A(n3845), .Y(n3798) );
  CLKBUFX3 U2851 ( .A(n3845), .Y(n3799) );
  CLKBUFX3 U2852 ( .A(n3845), .Y(n3800) );
  CLKBUFX3 U2853 ( .A(n3845), .Y(n3801) );
  CLKBUFX3 U2854 ( .A(n3844), .Y(n3802) );
  CLKBUFX3 U2855 ( .A(n3844), .Y(n3803) );
  CLKBUFX3 U2856 ( .A(n3844), .Y(n3804) );
  CLKBUFX3 U2857 ( .A(n3844), .Y(n3805) );
  CLKBUFX3 U2858 ( .A(n3843), .Y(n3806) );
  CLKBUFX3 U2859 ( .A(n3843), .Y(n3807) );
  CLKBUFX3 U2860 ( .A(n3843), .Y(n3808) );
  CLKBUFX3 U2861 ( .A(n3843), .Y(n3809) );
  CLKBUFX3 U2862 ( .A(n3842), .Y(n3810) );
  CLKBUFX3 U2863 ( .A(n3842), .Y(n3811) );
  CLKBUFX3 U2864 ( .A(n3842), .Y(n3812) );
  CLKBUFX3 U2865 ( .A(n3842), .Y(n3813) );
  CLKBUFX3 U2866 ( .A(n3841), .Y(n3814) );
  CLKBUFX3 U2867 ( .A(n3841), .Y(n3815) );
  CLKBUFX3 U2868 ( .A(n3841), .Y(n3816) );
  CLKBUFX3 U2869 ( .A(n3841), .Y(n3817) );
  CLKBUFX3 U2870 ( .A(n3840), .Y(n3818) );
  CLKBUFX3 U2871 ( .A(n3840), .Y(n3819) );
  CLKBUFX3 U2872 ( .A(n3840), .Y(n3820) );
  CLKBUFX3 U2873 ( .A(n3840), .Y(n3821) );
  CLKBUFX3 U2874 ( .A(n3839), .Y(n3822) );
  CLKBUFX3 U2875 ( .A(n3839), .Y(n3823) );
  CLKBUFX3 U2876 ( .A(n3839), .Y(n3824) );
  CLKBUFX3 U2877 ( .A(n3839), .Y(n3825) );
  CLKBUFX3 U2878 ( .A(n3733), .Y(n3826) );
  CLKBUFX3 U2879 ( .A(n3733), .Y(n3827) );
  CLKBUFX3 U2880 ( .A(n3845), .Y(n3828) );
  CLKBUFX3 U2881 ( .A(n3843), .Y(n3829) );
  CLKBUFX3 U2882 ( .A(n4140), .Y(n3659) );
  CLKBUFX3 U2883 ( .A(n351), .Y(n3901) );
  CLKBUFX3 U2884 ( .A(n351), .Y(n3902) );
  INVX3 U2885 ( .A(n3870), .Y(n3868) );
  INVX3 U2886 ( .A(mem_write), .Y(n3867) );
  INVX3 U2887 ( .A(n3870), .Y(n3866) );
  INVX3 U2888 ( .A(n3870), .Y(n3865) );
  INVX3 U2889 ( .A(n3870), .Y(n3864) );
  INVX3 U2890 ( .A(n3870), .Y(n3863) );
  INVX3 U2891 ( .A(mem_write), .Y(n3862) );
  INVX3 U2892 ( .A(n3870), .Y(n3869) );
  CLKBUFX3 U2893 ( .A(n351), .Y(n3900) );
  CLKBUFX3 U2894 ( .A(n351), .Y(n3899) );
  CLKBUFX3 U2895 ( .A(n351), .Y(n3898) );
  CLKBUFX3 U2896 ( .A(n351), .Y(n3896) );
  CLKBUFX3 U2897 ( .A(n351), .Y(n3897) );
  CLKBUFX3 U2898 ( .A(n3930), .Y(n3929) );
  CLKBUFX3 U2899 ( .A(n4098), .Y(n4097) );
  CLKBUFX3 U2900 ( .A(n4042), .Y(n4041) );
  CLKBUFX3 U2901 ( .A(n3986), .Y(n3985) );
  CLKINVX1 U2902 ( .A(n347), .Y(n3957) );
  CLKINVX1 U2903 ( .A(n347), .Y(n3958) );
  CLKBUFX3 U2904 ( .A(n3838), .Y(n3830) );
  CLKBUFX3 U2905 ( .A(n3838), .Y(n3831) );
  CLKBUFX3 U2906 ( .A(n3838), .Y(n3832) );
  CLKBUFX3 U2907 ( .A(n3838), .Y(n3833) );
  CLKBUFX3 U2908 ( .A(n3861), .Y(n3834) );
  CLKBUFX3 U2909 ( .A(n3861), .Y(n3835) );
  CLKBUFX3 U2910 ( .A(n3730), .Y(n3836) );
  CLKBUFX3 U2911 ( .A(n3844), .Y(n3837) );
  CLKBUFX3 U2912 ( .A(n3861), .Y(n3860) );
  CLKBUFX3 U2913 ( .A(n3861), .Y(n3859) );
  CLKBUFX3 U2914 ( .A(n3729), .Y(n3858) );
  CLKBUFX3 U2915 ( .A(n3730), .Y(n3857) );
  CLKBUFX3 U2916 ( .A(n3730), .Y(n3856) );
  CLKBUFX3 U2917 ( .A(n3730), .Y(n3855) );
  CLKBUFX3 U2918 ( .A(n3731), .Y(n3854) );
  CLKBUFX3 U2919 ( .A(n3732), .Y(n3853) );
  CLKBUFX3 U2920 ( .A(n3731), .Y(n3852) );
  CLKBUFX3 U2921 ( .A(n3729), .Y(n3851) );
  CLKBUFX3 U2922 ( .A(n3731), .Y(n3850) );
  CLKBUFX3 U2923 ( .A(n3731), .Y(n3849) );
  CLKBUFX3 U2924 ( .A(n3732), .Y(n3848) );
  CLKBUFX3 U2925 ( .A(n3732), .Y(n3847) );
  CLKBUFX3 U2926 ( .A(n3733), .Y(n3846) );
  CLKBUFX3 U2927 ( .A(n3729), .Y(n3845) );
  CLKBUFX3 U2928 ( .A(n3730), .Y(n3844) );
  CLKBUFX3 U2929 ( .A(n3851), .Y(n3843) );
  CLKBUFX3 U2930 ( .A(n3858), .Y(n3842) );
  CLKBUFX3 U2931 ( .A(n3733), .Y(n3841) );
  CLKBUFX3 U2932 ( .A(n3861), .Y(n3840) );
  CLKBUFX3 U2933 ( .A(n3733), .Y(n3839) );
  CLKINVX1 U2934 ( .A(n533), .Y(n4144) );
  NOR2X1 U2935 ( .A(mem_read), .B(mem_write), .Y(n536) );
  CLKBUFX3 U2936 ( .A(n366), .Y(n3885) );
  CLKBUFX3 U2937 ( .A(n366), .Y(n3886) );
  CLKBUFX3 U2938 ( .A(n351), .Y(n3895) );
  CLKBUFX3 U2939 ( .A(n351), .Y(n3894) );
  CLKBUFX3 U2940 ( .A(n3873), .Y(mem_write) );
  CLKBUFX3 U2941 ( .A(n3873), .Y(n3870) );
  CLKBUFX3 U2942 ( .A(n3873), .Y(n3872) );
  CLKBUFX3 U2943 ( .A(n17), .Y(n4127) );
  CLKBUFX3 U2944 ( .A(n17), .Y(n4128) );
  CLKBUFX3 U2945 ( .A(n351), .Y(n3893) );
  CLKINVX1 U2946 ( .A(n349), .Y(n3930) );
  CLKINVX1 U2947 ( .A(n208), .Y(n4098) );
  CLKINVX1 U2948 ( .A(n341), .Y(n4042) );
  CLKINVX1 U2949 ( .A(n345), .Y(n3986) );
  CLKINVX1 U2950 ( .A(n177), .Y(n4126) );
  CLKINVX1 U2951 ( .A(n177), .Y(n4125) );
  CLKINVX1 U2952 ( .A(n338), .Y(n4069) );
  CLKINVX1 U2953 ( .A(n338), .Y(n4070) );
  CLKINVX1 U2954 ( .A(n343), .Y(n4013) );
  CLKINVX1 U2955 ( .A(n343), .Y(n4014) );
  CLKBUFX3 U2956 ( .A(n3729), .Y(n3861) );
  CLKBUFX3 U2957 ( .A(n3729), .Y(n3838) );
  OAI31XL U2958 ( .A0(n3341), .A1(n4146), .A2(n3314), .B0(n430), .Y(n355) );
  OA21X2 U2959 ( .A0(n362), .A1(n4145), .B0(n361), .Y(n206) );
  OAI221XL U2960 ( .A0(n4133), .A1(n3255), .B0(n4131), .B1(n3193), .C0(n116), 
        .Y(proc_rdata[1]) );
  OA22X1 U2961 ( .A0(n4130), .A1(n3279), .B0(n4127), .B1(n3239), .Y(n116) );
  OAI221XL U2962 ( .A0(n4133), .A1(n3256), .B0(n4131), .B1(n3194), .C0(n61), 
        .Y(proc_rdata[2]) );
  OA22X1 U2963 ( .A0(n4129), .A1(n3280), .B0(n4128), .B1(n3242), .Y(n61) );
  OAI221XL U2964 ( .A0(n4134), .A1(n3257), .B0(n4131), .B1(n3195), .C0(n46), 
        .Y(proc_rdata[3]) );
  OA22X1 U2965 ( .A0(n4130), .A1(n3281), .B0(n4128), .B1(n3240), .Y(n46) );
  OAI221XL U2966 ( .A0(n4133), .A1(n3258), .B0(n4131), .B1(n3196), .C0(n41), 
        .Y(proc_rdata[4]) );
  OA22X1 U2967 ( .A0(n4130), .A1(n3282), .B0(n4127), .B1(n3243), .Y(n41) );
  OAI221XL U2968 ( .A0(n4134), .A1(n3259), .B0(n4131), .B1(n3197), .C0(n36), 
        .Y(proc_rdata[5]) );
  OA22X1 U2969 ( .A0(n4130), .A1(n3283), .B0(n4128), .B1(n3235), .Y(n36) );
  OAI221XL U2970 ( .A0(n4133), .A1(n3260), .B0(n4131), .B1(n3198), .C0(n31), 
        .Y(proc_rdata[6]) );
  OA22X1 U2971 ( .A0(n4130), .A1(n3284), .B0(n4127), .B1(n3244), .Y(n31) );
  OAI221XL U2972 ( .A0(n4134), .A1(n3261), .B0(n4131), .B1(n3206), .C0(n26), 
        .Y(proc_rdata[7]) );
  OA22X1 U2973 ( .A0(n4130), .A1(n3285), .B0(n4128), .B1(n3237), .Y(n26) );
  OAI221XL U2974 ( .A0(n4133), .A1(n3262), .B0(n4131), .B1(n3207), .C0(n21), 
        .Y(proc_rdata[8]) );
  OA22X1 U2975 ( .A0(n4130), .A1(n3286), .B0(n4127), .B1(n3236), .Y(n21) );
  OAI221XL U2976 ( .A0(n10), .A1(n3263), .B0(n4131), .B1(n3208), .C0(n14), .Y(
        proc_rdata[9]) );
  OA22X1 U2977 ( .A0(n4130), .A1(n3287), .B0(n4128), .B1(n3238), .Y(n14) );
  OAI221XL U2978 ( .A0(n4133), .A1(n3271), .B0(n4132), .B1(n3216), .C0(n131), 
        .Y(proc_rdata[17]) );
  OA22X1 U2979 ( .A0(n4130), .A1(n3230), .B0(n4127), .B1(n3301), .Y(n131) );
  OAI221XL U2980 ( .A0(n4133), .A1(n3272), .B0(n4131), .B1(n3217), .C0(n126), 
        .Y(proc_rdata[18]) );
  OA22X1 U2981 ( .A0(n4130), .A1(n3231), .B0(n4127), .B1(n3302), .Y(n126) );
  OAI221XL U2982 ( .A0(n4133), .A1(n3273), .B0(n4132), .B1(n3218), .C0(n121), 
        .Y(proc_rdata[19]) );
  OA22X1 U2983 ( .A0(n4130), .A1(n3232), .B0(n4127), .B1(n3309), .Y(n121) );
  OAI221XL U2984 ( .A0(n4133), .A1(n3274), .B0(n4131), .B1(n3219), .C0(n111), 
        .Y(proc_rdata[20]) );
  OA22X1 U2985 ( .A0(n4129), .A1(n3233), .B0(n4128), .B1(n3303), .Y(n111) );
  OAI221XL U2986 ( .A0(n4133), .A1(n3275), .B0(n4132), .B1(n3220), .C0(n106), 
        .Y(proc_rdata[21]) );
  OA22X1 U2987 ( .A0(n4129), .A1(n3234), .B0(n4128), .B1(n3304), .Y(n106) );
  OAI221XL U2988 ( .A0(n4133), .A1(n3276), .B0(n4131), .B1(n3221), .C0(n101), 
        .Y(proc_rdata[22]) );
  OA22X1 U2989 ( .A0(n4129), .A1(n3223), .B0(n4128), .B1(n3305), .Y(n101) );
  OAI221XL U2990 ( .A0(n4133), .A1(n3277), .B0(n12), .B1(n3222), .C0(n96), .Y(
        proc_rdata[23]) );
  OA22X1 U2991 ( .A0(n4129), .A1(n3354), .B0(n4128), .B1(n3306), .Y(n96) );
  OAI221XL U2992 ( .A0(n4133), .A1(n3246), .B0(n4131), .B1(n3199), .C0(n91), 
        .Y(proc_rdata[24]) );
  OA22X1 U2993 ( .A0(n4129), .A1(n3357), .B0(n4128), .B1(n3289), .Y(n91) );
  OAI221XL U2994 ( .A0(n4133), .A1(n3247), .B0(n4132), .B1(n3200), .C0(n86), 
        .Y(proc_rdata[25]) );
  OA22X1 U2995 ( .A0(n4129), .A1(n3360), .B0(n4128), .B1(n3290), .Y(n86) );
  OAI221XL U2996 ( .A0(n4133), .A1(n3248), .B0(n4131), .B1(n3201), .C0(n81), 
        .Y(proc_rdata[26]) );
  OA22X1 U2997 ( .A0(n4129), .A1(n3363), .B0(n4128), .B1(n3291), .Y(n81) );
  OAI221XL U2998 ( .A0(n4133), .A1(n3249), .B0(n4132), .B1(n3202), .C0(n76), 
        .Y(proc_rdata[27]) );
  OA22X1 U2999 ( .A0(n4129), .A1(n3366), .B0(n4128), .B1(n3292), .Y(n76) );
  OAI221XL U3000 ( .A0(n4133), .A1(n3250), .B0(n4131), .B1(n3203), .C0(n71), 
        .Y(proc_rdata[28]) );
  OA22X1 U3001 ( .A0(n4129), .A1(n3369), .B0(n4128), .B1(n3293), .Y(n71) );
  OAI221XL U3002 ( .A0(n4134), .A1(n3251), .B0(n4131), .B1(n3204), .C0(n66), 
        .Y(proc_rdata[29]) );
  OA22X1 U3003 ( .A0(n4129), .A1(n3372), .B0(n4128), .B1(n3294), .Y(n66) );
  OAI221XL U3004 ( .A0(n4133), .A1(n3252), .B0(n4131), .B1(n3205), .C0(n56), 
        .Y(proc_rdata[30]) );
  OA22X1 U3005 ( .A0(n4129), .A1(n3375), .B0(n4128), .B1(n3295), .Y(n56) );
  OAI221XL U3006 ( .A0(n4134), .A1(n3253), .B0(n4131), .B1(n3191), .C0(n51), 
        .Y(proc_rdata[31]) );
  OA22X1 U3007 ( .A0(n4130), .A1(n3378), .B0(n4127), .B1(n3296), .Y(n51) );
  OAI221XL U3008 ( .A0(n4134), .A1(n3254), .B0(n4132), .B1(n3192), .C0(n171), 
        .Y(proc_rdata[0]) );
  OA22X1 U3009 ( .A0(n4129), .A1(n3278), .B0(n4127), .B1(n3190), .Y(n171) );
  OAI221XL U3010 ( .A0(n4134), .A1(n3264), .B0(n4132), .B1(n3209), .C0(n166), 
        .Y(proc_rdata[10]) );
  OA22X1 U3011 ( .A0(n4130), .A1(n3288), .B0(n4127), .B1(n3241), .Y(n166) );
  OAI221XL U3012 ( .A0(n4134), .A1(n3265), .B0(n4132), .B1(n3210), .C0(n161), 
        .Y(proc_rdata[11]) );
  OA22X1 U3013 ( .A0(n4129), .A1(n3224), .B0(n4127), .B1(n3297), .Y(n161) );
  OAI221XL U3014 ( .A0(n4134), .A1(n3266), .B0(n4132), .B1(n3211), .C0(n156), 
        .Y(proc_rdata[12]) );
  OA22X1 U3015 ( .A0(n4130), .A1(n3225), .B0(n4127), .B1(n3307), .Y(n156) );
  OAI221XL U3016 ( .A0(n4134), .A1(n3267), .B0(n4132), .B1(n3212), .C0(n151), 
        .Y(proc_rdata[13]) );
  OA22X1 U3017 ( .A0(n4129), .A1(n3226), .B0(n4127), .B1(n3308), .Y(n151) );
  OAI221XL U3018 ( .A0(n4134), .A1(n3268), .B0(n4132), .B1(n3213), .C0(n146), 
        .Y(proc_rdata[14]) );
  OA22X1 U3019 ( .A0(n4130), .A1(n3227), .B0(n4127), .B1(n3298), .Y(n146) );
  OAI221XL U3020 ( .A0(n4134), .A1(n3269), .B0(n4132), .B1(n3214), .C0(n141), 
        .Y(proc_rdata[15]) );
  OA22X1 U3021 ( .A0(n4129), .A1(n3228), .B0(n4127), .B1(n3299), .Y(n141) );
  OAI221XL U3022 ( .A0(n4134), .A1(n3270), .B0(n4132), .B1(n3215), .C0(n136), 
        .Y(proc_rdata[16]) );
  OA22X1 U3023 ( .A0(n4130), .A1(n3229), .B0(n4127), .B1(n3300), .Y(n136) );
  NAND3X2 U3024 ( .A(n4146), .B(n3314), .C(n4143), .Y(n366) );
  CLKINVX1 U3025 ( .A(n361), .Y(n4143) );
  CLKINVX1 U3026 ( .A(N34), .Y(n4145) );
  CLKBUFX3 U3027 ( .A(n358), .Y(n3888) );
  CLKBUFX3 U3028 ( .A(n358), .Y(n3889) );
  CLKBUFX3 U3029 ( .A(n353), .Y(n3891) );
  CLKBUFX3 U3030 ( .A(n467), .Y(n3874) );
  CLKBUFX3 U3031 ( .A(n467), .Y(n3875) );
  CLKBUFX3 U3032 ( .A(n12), .Y(n4131) );
  CLKBUFX3 U3033 ( .A(n10), .Y(n4133) );
  CLKBUFX3 U3034 ( .A(n15), .Y(n4129) );
  NOR2X1 U3035 ( .A(n3192), .B(n3864), .Y(mem_wdata[64]) );
  NOR2X1 U3036 ( .A(n3193), .B(n3864), .Y(mem_wdata[65]) );
  NOR2X1 U3037 ( .A(n3194), .B(n3864), .Y(mem_wdata[66]) );
  NOR2X1 U3038 ( .A(n3195), .B(n3864), .Y(mem_wdata[67]) );
  NOR2X1 U3039 ( .A(n3196), .B(n3863), .Y(mem_wdata[68]) );
  NOR2X1 U3040 ( .A(n3197), .B(n3863), .Y(mem_wdata[69]) );
  NOR2X1 U3041 ( .A(n3198), .B(n3863), .Y(mem_wdata[70]) );
  NOR2X1 U3042 ( .A(n3206), .B(n3863), .Y(mem_wdata[71]) );
  NOR2X1 U3043 ( .A(n3207), .B(n3863), .Y(mem_wdata[72]) );
  NOR2X1 U3044 ( .A(n3208), .B(n3863), .Y(mem_wdata[73]) );
  NOR2X1 U3045 ( .A(n3209), .B(n3863), .Y(mem_wdata[74]) );
  NOR2X1 U3046 ( .A(n3210), .B(n3863), .Y(mem_wdata[75]) );
  NOR2X1 U3047 ( .A(n3211), .B(n3863), .Y(mem_wdata[76]) );
  NOR2X1 U3048 ( .A(n3212), .B(n3863), .Y(mem_wdata[77]) );
  NOR2X1 U3049 ( .A(n3213), .B(n3863), .Y(mem_wdata[78]) );
  NOR2X1 U3050 ( .A(n3214), .B(n3864), .Y(mem_wdata[79]) );
  NOR2X1 U3051 ( .A(n3215), .B(n3863), .Y(mem_wdata[80]) );
  NOR2X1 U3052 ( .A(n3216), .B(n3864), .Y(mem_wdata[81]) );
  NOR2X1 U3053 ( .A(n3217), .B(n3863), .Y(mem_wdata[82]) );
  NOR2X1 U3054 ( .A(n3218), .B(n3864), .Y(mem_wdata[83]) );
  NOR2X1 U3055 ( .A(n3219), .B(n3863), .Y(mem_wdata[84]) );
  NOR2X1 U3056 ( .A(n3220), .B(n3865), .Y(mem_wdata[85]) );
  NOR2X1 U3057 ( .A(n3221), .B(n3869), .Y(mem_wdata[86]) );
  NOR2X1 U3058 ( .A(n3222), .B(n3867), .Y(mem_wdata[87]) );
  NOR2X1 U3059 ( .A(n3199), .B(n3862), .Y(mem_wdata[88]) );
  NOR2X1 U3060 ( .A(n3200), .B(n3864), .Y(mem_wdata[89]) );
  NOR2X1 U3061 ( .A(n3201), .B(n3862), .Y(mem_wdata[90]) );
  NOR2X1 U3062 ( .A(n3202), .B(n3862), .Y(mem_wdata[91]) );
  NOR2X1 U3063 ( .A(n3203), .B(n3862), .Y(mem_wdata[92]) );
  NOR2X1 U3064 ( .A(n3204), .B(n3862), .Y(mem_wdata[93]) );
  NOR2X1 U3065 ( .A(n3205), .B(n3862), .Y(mem_wdata[94]) );
  NOR2X1 U3066 ( .A(n3191), .B(n3862), .Y(mem_wdata[95]) );
  NOR2X1 U3067 ( .A(n3254), .B(n3867), .Y(mem_wdata[32]) );
  NOR2X1 U3068 ( .A(n3255), .B(n3867), .Y(mem_wdata[33]) );
  NOR2X1 U3069 ( .A(n3256), .B(n3867), .Y(mem_wdata[34]) );
  NOR2X1 U3070 ( .A(n3257), .B(n3866), .Y(mem_wdata[35]) );
  NOR2X1 U3071 ( .A(n3258), .B(n3866), .Y(mem_wdata[36]) );
  NOR2X1 U3072 ( .A(n3259), .B(n3866), .Y(mem_wdata[37]) );
  NOR2X1 U3073 ( .A(n3260), .B(n3866), .Y(mem_wdata[38]) );
  NOR2X1 U3074 ( .A(n3261), .B(n3866), .Y(mem_wdata[39]) );
  NOR2X1 U3075 ( .A(n3262), .B(n3866), .Y(mem_wdata[40]) );
  NOR2X1 U3076 ( .A(n3263), .B(n3866), .Y(mem_wdata[41]) );
  NOR2X1 U3077 ( .A(n3264), .B(n3866), .Y(mem_wdata[42]) );
  NOR2X1 U3078 ( .A(n3265), .B(n3866), .Y(mem_wdata[43]) );
  NOR2X1 U3079 ( .A(n3266), .B(n3866), .Y(mem_wdata[44]) );
  NOR2X1 U3080 ( .A(n3267), .B(n3866), .Y(mem_wdata[45]) );
  NOR2X1 U3081 ( .A(n3268), .B(n3865), .Y(mem_wdata[46]) );
  NOR2X1 U3082 ( .A(n3269), .B(n3865), .Y(mem_wdata[47]) );
  NOR2X1 U3083 ( .A(n3270), .B(n3865), .Y(mem_wdata[48]) );
  NOR2X1 U3084 ( .A(n3271), .B(n3865), .Y(mem_wdata[49]) );
  NOR2X1 U3085 ( .A(n3272), .B(n3865), .Y(mem_wdata[50]) );
  NOR2X1 U3086 ( .A(n3273), .B(n3865), .Y(mem_wdata[51]) );
  NOR2X1 U3087 ( .A(n3274), .B(n3865), .Y(mem_wdata[52]) );
  NOR2X1 U3088 ( .A(n3275), .B(n3865), .Y(mem_wdata[53]) );
  NOR2X1 U3089 ( .A(n3276), .B(n3865), .Y(mem_wdata[54]) );
  NOR2X1 U3090 ( .A(n3277), .B(n3865), .Y(mem_wdata[55]) );
  NOR2X1 U3091 ( .A(n3246), .B(n3865), .Y(mem_wdata[56]) );
  NOR2X1 U3092 ( .A(n3247), .B(n3864), .Y(mem_wdata[57]) );
  NOR2X1 U3093 ( .A(n3248), .B(n3864), .Y(mem_wdata[58]) );
  NOR2X1 U3094 ( .A(n3249), .B(n3864), .Y(mem_wdata[59]) );
  NOR2X1 U3095 ( .A(n3250), .B(n3864), .Y(mem_wdata[60]) );
  NOR2X1 U3096 ( .A(n3251), .B(n3864), .Y(mem_wdata[61]) );
  NOR2X1 U3097 ( .A(n3252), .B(n3864), .Y(mem_wdata[62]) );
  NOR2X1 U3098 ( .A(n3253), .B(n3864), .Y(mem_wdata[63]) );
  NOR2X1 U3099 ( .A(n3190), .B(n3869), .Y(mem_wdata[0]) );
  NOR2X1 U3100 ( .A(n3239), .B(n3868), .Y(mem_wdata[1]) );
  NOR2X1 U3101 ( .A(n3242), .B(n3867), .Y(mem_wdata[2]) );
  NOR2X1 U3102 ( .A(n3240), .B(n3866), .Y(mem_wdata[3]) );
  NOR2X1 U3103 ( .A(n3243), .B(n3865), .Y(mem_wdata[4]) );
  NOR2X1 U3104 ( .A(n3235), .B(n3864), .Y(mem_wdata[5]) );
  NOR2X1 U3105 ( .A(n3244), .B(n3863), .Y(mem_wdata[6]) );
  NOR2X1 U3106 ( .A(n3237), .B(n3863), .Y(mem_wdata[7]) );
  NOR2X1 U3107 ( .A(n3236), .B(n3862), .Y(mem_wdata[8]) );
  NOR2X1 U3108 ( .A(n3238), .B(n3862), .Y(mem_wdata[9]) );
  NOR2X1 U3109 ( .A(n3241), .B(n3867), .Y(mem_wdata[10]) );
  NOR2X1 U3110 ( .A(n3297), .B(n3869), .Y(mem_wdata[11]) );
  NOR2X1 U3111 ( .A(n3307), .B(n3869), .Y(mem_wdata[12]) );
  NOR2X1 U3112 ( .A(n3308), .B(n3868), .Y(mem_wdata[13]) );
  NOR2X1 U3113 ( .A(n3298), .B(n3868), .Y(mem_wdata[14]) );
  NOR2X1 U3114 ( .A(n3299), .B(n3868), .Y(mem_wdata[15]) );
  NOR2X1 U3115 ( .A(n3300), .B(n3868), .Y(mem_wdata[16]) );
  NOR2X1 U3116 ( .A(n3301), .B(n3868), .Y(mem_wdata[17]) );
  NOR2X1 U3117 ( .A(n3302), .B(n3868), .Y(mem_wdata[18]) );
  NOR2X1 U3118 ( .A(n3309), .B(n3868), .Y(mem_wdata[19]) );
  NOR2X1 U3119 ( .A(n3303), .B(n3868), .Y(mem_wdata[20]) );
  NOR2X1 U3120 ( .A(n3304), .B(n3868), .Y(mem_wdata[21]) );
  NOR2X1 U3121 ( .A(n3305), .B(n3868), .Y(mem_wdata[22]) );
  NOR2X1 U3122 ( .A(n3306), .B(n3868), .Y(mem_wdata[23]) );
  NOR2X1 U3123 ( .A(n3289), .B(n3867), .Y(mem_wdata[24]) );
  NOR2X1 U3124 ( .A(n3290), .B(n3867), .Y(mem_wdata[25]) );
  NOR2X1 U3125 ( .A(n3291), .B(n3867), .Y(mem_wdata[26]) );
  NOR2X1 U3126 ( .A(n3292), .B(n3867), .Y(mem_wdata[27]) );
  NOR2X1 U3127 ( .A(n3293), .B(n3867), .Y(mem_wdata[28]) );
  NOR2X1 U3128 ( .A(n3294), .B(n3867), .Y(mem_wdata[29]) );
  NOR2X1 U3129 ( .A(n3295), .B(n3867), .Y(mem_wdata[30]) );
  NOR2X1 U3130 ( .A(n3296), .B(n3867), .Y(mem_wdata[31]) );
  NOR2X1 U3131 ( .A(n3278), .B(n3862), .Y(mem_wdata[96]) );
  NOR2X1 U3132 ( .A(n3279), .B(n3862), .Y(mem_wdata[97]) );
  NOR2X1 U3133 ( .A(n3280), .B(n3862), .Y(mem_wdata[98]) );
  NOR2X1 U3134 ( .A(n3281), .B(n3862), .Y(mem_wdata[99]) );
  NOR2X1 U3135 ( .A(n3282), .B(n3866), .Y(mem_wdata[100]) );
  NOR2X1 U3136 ( .A(n3283), .B(n3868), .Y(mem_wdata[101]) );
  NOR2X1 U3137 ( .A(n3284), .B(n3868), .Y(mem_wdata[102]) );
  NOR2X1 U3138 ( .A(n3285), .B(n3867), .Y(mem_wdata[103]) );
  NOR2X1 U3139 ( .A(n3286), .B(n3865), .Y(mem_wdata[104]) );
  NOR2X1 U3140 ( .A(n3287), .B(n3869), .Y(mem_wdata[105]) );
  NOR2X1 U3141 ( .A(n3288), .B(n3866), .Y(mem_wdata[106]) );
  NOR2X1 U3142 ( .A(n3224), .B(n3865), .Y(mem_wdata[107]) );
  NOR2X1 U3143 ( .A(n3225), .B(n3868), .Y(mem_wdata[108]) );
  NOR2X1 U3144 ( .A(n3226), .B(n3867), .Y(mem_wdata[109]) );
  NOR2X1 U3145 ( .A(n3227), .B(n3865), .Y(mem_wdata[110]) );
  NOR2X1 U3146 ( .A(n3228), .B(n3869), .Y(mem_wdata[111]) );
  NOR2X1 U3147 ( .A(n3229), .B(n3866), .Y(mem_wdata[112]) );
  NOR2X1 U3148 ( .A(n3230), .B(n3868), .Y(mem_wdata[113]) );
  NOR2X1 U3149 ( .A(n3231), .B(n3867), .Y(mem_wdata[114]) );
  NOR2X1 U3150 ( .A(n3232), .B(n3865), .Y(mem_wdata[115]) );
  NOR2X1 U3151 ( .A(n3233), .B(n3869), .Y(mem_wdata[116]) );
  NOR2X1 U3152 ( .A(n3234), .B(n3866), .Y(mem_wdata[117]) );
  NOR2X1 U3153 ( .A(n3223), .B(n3869), .Y(mem_wdata[118]) );
  NOR2X1 U3154 ( .A(n3354), .B(n3869), .Y(mem_wdata[119]) );
  NOR2X1 U3155 ( .A(n3357), .B(n3869), .Y(mem_wdata[120]) );
  NOR2X1 U3156 ( .A(n3360), .B(n3869), .Y(mem_wdata[121]) );
  NOR2X1 U3157 ( .A(n3363), .B(n3869), .Y(mem_wdata[122]) );
  NOR2X1 U3158 ( .A(n3366), .B(n3869), .Y(mem_wdata[123]) );
  NOR2X1 U3159 ( .A(n3369), .B(n3869), .Y(mem_wdata[124]) );
  NOR2X1 U3160 ( .A(n3372), .B(n3869), .Y(mem_wdata[125]) );
  NOR2X1 U3161 ( .A(n3375), .B(n3869), .Y(mem_wdata[126]) );
  NOR2X1 U3162 ( .A(n3378), .B(n3869), .Y(mem_wdata[127]) );
  NOR2X1 U3163 ( .A(n536), .B(n4139), .Y(mem_addr[1]) );
  NOR2X1 U3164 ( .A(n536), .B(n4137), .Y(mem_addr[2]) );
  CLKBUFX3 U3165 ( .A(n15), .Y(n4130) );
  CLKBUFX3 U3166 ( .A(n4142), .Y(n3729) );
  CLKBUFX3 U3167 ( .A(n4142), .Y(n3730) );
  CLKBUFX3 U3168 ( .A(n4142), .Y(n3731) );
  CLKBUFX3 U3169 ( .A(n4142), .Y(n3732) );
  CLKBUFX3 U3170 ( .A(n4142), .Y(n3733) );
  AOI21X2 U3171 ( .A0(mem_rdata[24]), .A1(n3899), .B0(n415), .Y(n234) );
  OAI22XL U3172 ( .A0(n3887), .A1(n4154), .B0(n3289), .B1(n3883), .Y(n415) );
  AOI21X2 U3173 ( .A0(mem_rdata[25]), .A1(n3899), .B0(n417), .Y(n235) );
  OAI22XL U3174 ( .A0(n3887), .A1(n4153), .B0(n3290), .B1(n3882), .Y(n417) );
  AOI21X2 U3175 ( .A0(mem_rdata[26]), .A1(n3899), .B0(n419), .Y(n236) );
  OAI22XL U3176 ( .A0(n3887), .A1(n4152), .B0(n3291), .B1(n3882), .Y(n419) );
  AOI21X2 U3177 ( .A0(mem_rdata[27]), .A1(n3899), .B0(n421), .Y(n237) );
  OAI22XL U3178 ( .A0(n3887), .A1(n4151), .B0(n3292), .B1(n3882), .Y(n421) );
  AOI21X2 U3179 ( .A0(mem_rdata[28]), .A1(n3899), .B0(n423), .Y(n238) );
  OAI22XL U3180 ( .A0(n3887), .A1(n4150), .B0(n3293), .B1(n3882), .Y(n423) );
  AOI21X2 U3181 ( .A0(mem_rdata[29]), .A1(n3899), .B0(n425), .Y(n239) );
  OAI22XL U3182 ( .A0(n3887), .A1(n4149), .B0(n3294), .B1(n3882), .Y(n425) );
  AOI21X2 U3183 ( .A0(mem_rdata[30]), .A1(n3899), .B0(n427), .Y(n240) );
  OAI22XL U3184 ( .A0(n4148), .A1(n3887), .B0(n3295), .B1(n3882), .Y(n427) );
  OAI22XL U3185 ( .A0(n4147), .A1(n3887), .B0(n3296), .B1(n3883), .Y(n428) );
  AOI21X2 U3186 ( .A0(mem_rdata[56]), .A1(n3893), .B0(n458), .Y(n266) );
  OAI22XL U3187 ( .A0(n4154), .A1(n3881), .B0(n3246), .B1(n3878), .Y(n458) );
  AOI21X2 U3188 ( .A0(mem_rdata[57]), .A1(n3893), .B0(n459), .Y(n267) );
  OAI22XL U3189 ( .A0(n4153), .A1(n3881), .B0(n3247), .B1(n3877), .Y(n459) );
  AOI21X2 U3190 ( .A0(mem_rdata[58]), .A1(n3893), .B0(n460), .Y(n268) );
  OAI22XL U3191 ( .A0(n4152), .A1(n3881), .B0(n3248), .B1(n434), .Y(n460) );
  AOI21X2 U3192 ( .A0(mem_rdata[59]), .A1(n3893), .B0(n461), .Y(n269) );
  OAI22XL U3193 ( .A0(n4151), .A1(n3881), .B0(n3249), .B1(n3878), .Y(n461) );
  AOI21X2 U3194 ( .A0(mem_rdata[60]), .A1(n3893), .B0(n462), .Y(n270) );
  OAI22XL U3195 ( .A0(n4150), .A1(n3881), .B0(n3250), .B1(n3877), .Y(n462) );
  AOI21X2 U3196 ( .A0(mem_rdata[61]), .A1(n3893), .B0(n463), .Y(n271) );
  OAI22XL U3197 ( .A0(n4149), .A1(n3881), .B0(n3251), .B1(n3878), .Y(n463) );
  AOI21X2 U3198 ( .A0(mem_rdata[62]), .A1(n3893), .B0(n464), .Y(n272) );
  OAI22XL U3199 ( .A0(n4148), .A1(n3881), .B0(n3252), .B1(n3877), .Y(n464) );
  AOI21X2 U3200 ( .A0(mem_rdata[63]), .A1(n3893), .B0(n465), .Y(n273) );
  OAI22XL U3201 ( .A0(n4147), .A1(n3881), .B0(n3253), .B1(n434), .Y(n465) );
  AOI21X2 U3202 ( .A0(mem_rdata[88]), .A1(n3900), .B0(n492), .Y(n298) );
  OAI22XL U3203 ( .A0(n4154), .A1(n3876), .B0(n3199), .B1(n3087), .Y(n492) );
  AOI21X2 U3204 ( .A0(mem_rdata[89]), .A1(n3895), .B0(n493), .Y(n299) );
  OAI22XL U3205 ( .A0(n4153), .A1(n3876), .B0(n3200), .B1(n3087), .Y(n493) );
  AOI21X2 U3206 ( .A0(mem_rdata[90]), .A1(n3896), .B0(n494), .Y(n300) );
  OAI22XL U3207 ( .A0(n4152), .A1(n3876), .B0(n3201), .B1(n3087), .Y(n494) );
  AOI21X2 U3208 ( .A0(mem_rdata[91]), .A1(n3896), .B0(n495), .Y(n301) );
  OAI22XL U3209 ( .A0(n4151), .A1(n3876), .B0(n3202), .B1(n3087), .Y(n495) );
  AOI21X2 U3210 ( .A0(mem_rdata[92]), .A1(n3896), .B0(n496), .Y(n302) );
  OAI22XL U3211 ( .A0(n4150), .A1(n3876), .B0(n3203), .B1(n3087), .Y(n496) );
  AOI21X2 U3212 ( .A0(mem_rdata[93]), .A1(n3896), .B0(n497), .Y(n303) );
  OAI22XL U3213 ( .A0(n4149), .A1(n3876), .B0(n3204), .B1(n3087), .Y(n497) );
  AOI21X2 U3214 ( .A0(mem_rdata[94]), .A1(n3896), .B0(n498), .Y(n304) );
  OAI22XL U3215 ( .A0(n4148), .A1(n3876), .B0(n3205), .B1(n3087), .Y(n498) );
  AOI21X2 U3216 ( .A0(mem_rdata[95]), .A1(n3896), .B0(n499), .Y(n305) );
  OAI22XL U3217 ( .A0(n4147), .A1(n3876), .B0(n3191), .B1(n3087), .Y(n499) );
  AOI21X2 U3218 ( .A0(mem_rdata[118]), .A1(n3894), .B0(n522), .Y(n328) );
  OAI22XL U3219 ( .A0(n3892), .A1(n4156), .B0(n3223), .B1(n3075), .Y(n522) );
  AOI21X2 U3220 ( .A0(mem_rdata[119]), .A1(n3894), .B0(n523), .Y(n329) );
  OAI22XL U3221 ( .A0(n3892), .A1(n4155), .B0(n3354), .B1(n3075), .Y(n523) );
  AOI21X2 U3222 ( .A0(mem_rdata[120]), .A1(n3894), .B0(n524), .Y(n330) );
  OAI22XL U3223 ( .A0(n3892), .A1(n4154), .B0(n3357), .B1(n3075), .Y(n524) );
  AOI21X2 U3224 ( .A0(mem_rdata[121]), .A1(n3894), .B0(n525), .Y(n331) );
  OAI22XL U3225 ( .A0(n3892), .A1(n4153), .B0(n3360), .B1(n3075), .Y(n525) );
  AOI21X2 U3226 ( .A0(mem_rdata[122]), .A1(n3894), .B0(n526), .Y(n332) );
  AOI21X2 U3227 ( .A0(mem_rdata[123]), .A1(n3894), .B0(n527), .Y(n333) );
  OAI22XL U3228 ( .A0(n3892), .A1(n4151), .B0(n3366), .B1(n3075), .Y(n527) );
  AOI21X2 U3229 ( .A0(mem_rdata[124]), .A1(n3894), .B0(n528), .Y(n334) );
  OAI22XL U3230 ( .A0(n3892), .A1(n4150), .B0(n3369), .B1(n3075), .Y(n528) );
  AOI21X2 U3231 ( .A0(mem_rdata[125]), .A1(n3897), .B0(n529), .Y(n335) );
  OAI22XL U3232 ( .A0(n3892), .A1(n4149), .B0(n3372), .B1(n3075), .Y(n529) );
  MXI2X1 U3233 ( .A(n3625), .B(n3626), .S0(n3726), .Y(N57) );
  MXI2X1 U3234 ( .A(n3631), .B(n3632), .S0(n3727), .Y(N54) );
  MXI2X1 U3235 ( .A(n3633), .B(n3634), .S0(n3727), .Y(N53) );
  MXI2X1 U3236 ( .A(n3635), .B(n3636), .S0(n3727), .Y(N52) );
  MXI4X1 U3237 ( .A(\CACHE[0][135] ), .B(\CACHE[1][135] ), .C(\CACHE[2][135] ), 
        .D(\CACHE[3][135] ), .S0(n3683), .S1(n3689), .Y(n3635) );
  MXI4X1 U3238 ( .A(\CACHE[4][129] ), .B(\CACHE[5][129] ), .C(\CACHE[6][129] ), 
        .D(\CACHE[7][129] ), .S0(n3682), .S1(n3711), .Y(n3624) );
  MXI2X1 U3239 ( .A(n3629), .B(n3630), .S0(n3727), .Y(N55) );
  MXI2X1 U3240 ( .A(n3637), .B(n3638), .S0(n3727), .Y(N51) );
  MXI2X1 U3241 ( .A(n3639), .B(n3640), .S0(n3727), .Y(N50) );
  MXI2X1 U3242 ( .A(n3641), .B(n3642), .S0(n3727), .Y(N49) );
  MXI2X1 U3243 ( .A(n3643), .B(n3644), .S0(n3727), .Y(N48) );
  MXI2X1 U3244 ( .A(n3645), .B(n3646), .S0(n3727), .Y(N46) );
  MXI2X1 U3245 ( .A(n3647), .B(n3648), .S0(n3727), .Y(N45) );
  MXI2X1 U3246 ( .A(n3649), .B(n3650), .S0(n3728), .Y(N44) );
  MXI2X1 U3247 ( .A(n3653), .B(n3654), .S0(n3728), .Y(N38) );
  MXI4X1 U3248 ( .A(\CACHE[0][149] ), .B(\CACHE[1][149] ), .C(\CACHE[2][149] ), 
        .D(\CACHE[3][149] ), .S0(n3685), .S1(n3715), .Y(n3653) );
  MXI4X1 U3249 ( .A(\CACHE[4][149] ), .B(\CACHE[5][149] ), .C(\CACHE[6][149] ), 
        .D(\CACHE[7][149] ), .S0(n3685), .S1(n3715), .Y(n3654) );
  XOR2X1 U3250 ( .A(proc_addr[27]), .B(N37), .Y(n546) );
  XOR2X1 U3251 ( .A(proc_addr[21]), .B(N43), .Y(n554) );
  XOR2X1 U3252 ( .A(proc_addr[10]), .B(N54), .Y(n561) );
  XOR2X1 U3253 ( .A(proc_addr[12]), .B(N52), .Y(n568) );
  XOR2X1 U3254 ( .A(proc_addr[22]), .B(N42), .Y(n553) );
  XOR2X1 U3255 ( .A(proc_addr[29]), .B(N35), .Y(n560) );
  XOR2X1 U3256 ( .A(proc_addr[11]), .B(N53), .Y(n567) );
  XOR2X1 U3257 ( .A(proc_addr[24]), .B(N40), .Y(n552) );
  XOR2X1 U3258 ( .A(proc_addr[23]), .B(N41), .Y(n559) );
  XOR2X1 U3259 ( .A(proc_addr[7]), .B(N57), .Y(n566) );
  XNOR2X1 U3260 ( .A(N59), .B(proc_addr[5]), .Y(n550) );
  XOR2X1 U3261 ( .A(proc_addr[28]), .B(N36), .Y(n544) );
  XOR2X1 U3262 ( .A(proc_addr[17]), .B(N47), .Y(n545) );
  XNOR2X1 U3263 ( .A(N58), .B(proc_addr[6]), .Y(n549) );
  XNOR2X1 U3264 ( .A(N56), .B(proc_addr[8]), .Y(n548) );
  AOI21X2 U3265 ( .A0(mem_rdata[0]), .A1(n3901), .B0(n365), .Y(n209) );
  OAI22XL U3266 ( .A0(n3885), .A1(n4177), .B0(n3239), .B1(n3883), .Y(n369) );
  AOI21X2 U3267 ( .A0(mem_rdata[2]), .A1(n3901), .B0(n371), .Y(n212) );
  OAI22XL U3268 ( .A0(n3885), .A1(n4176), .B0(n3242), .B1(n3883), .Y(n371) );
  AOI21X2 U3269 ( .A0(mem_rdata[3]), .A1(n3901), .B0(n373), .Y(n213) );
  OAI22XL U3270 ( .A0(n3885), .A1(n4175), .B0(n3240), .B1(n3883), .Y(n373) );
  AOI21X2 U3271 ( .A0(mem_rdata[4]), .A1(n3901), .B0(n375), .Y(n214) );
  OAI22XL U3272 ( .A0(n3885), .A1(n4174), .B0(n3243), .B1(n3883), .Y(n375) );
  AOI21X2 U3273 ( .A0(mem_rdata[5]), .A1(n3901), .B0(n377), .Y(n215) );
  OAI22XL U3274 ( .A0(n3885), .A1(n4173), .B0(n3235), .B1(n3883), .Y(n377) );
  AOI21X2 U3275 ( .A0(mem_rdata[6]), .A1(n3901), .B0(n379), .Y(n216) );
  OAI22XL U3276 ( .A0(n3885), .A1(n4172), .B0(n3244), .B1(n3883), .Y(n379) );
  AOI21X2 U3277 ( .A0(mem_rdata[7]), .A1(n3900), .B0(n381), .Y(n217) );
  OAI22XL U3278 ( .A0(n3885), .A1(n4171), .B0(n3237), .B1(n3883), .Y(n381) );
  AOI21X2 U3279 ( .A0(mem_rdata[8]), .A1(n3900), .B0(n383), .Y(n218) );
  OAI22XL U3280 ( .A0(n3885), .A1(n4170), .B0(n3236), .B1(n3883), .Y(n383) );
  AOI21X2 U3281 ( .A0(mem_rdata[9]), .A1(n3900), .B0(n385), .Y(n219) );
  OAI22XL U3282 ( .A0(n3885), .A1(n4169), .B0(n3238), .B1(n3883), .Y(n385) );
  AOI21X2 U3283 ( .A0(mem_rdata[10]), .A1(n3900), .B0(n387), .Y(n220) );
  OAI22XL U3284 ( .A0(n3885), .A1(n4168), .B0(n3241), .B1(n3883), .Y(n387) );
  AOI21X2 U3285 ( .A0(mem_rdata[11]), .A1(n3900), .B0(n389), .Y(n221) );
  OAI22XL U3286 ( .A0(n3885), .A1(n4167), .B0(n3297), .B1(n3883), .Y(n389) );
  AOI21X2 U3287 ( .A0(mem_rdata[14]), .A1(n3900), .B0(n395), .Y(n224) );
  OAI22XL U3288 ( .A0(n3886), .A1(n4164), .B0(n3298), .B1(n3884), .Y(n395) );
  AOI21X2 U3289 ( .A0(mem_rdata[15]), .A1(n3900), .B0(n397), .Y(n225) );
  OAI22XL U3290 ( .A0(n3886), .A1(n4163), .B0(n3299), .B1(n3884), .Y(n397) );
  AOI21X2 U3291 ( .A0(mem_rdata[16]), .A1(n3900), .B0(n399), .Y(n226) );
  OAI22XL U3292 ( .A0(n3886), .A1(n4162), .B0(n3300), .B1(n3884), .Y(n399) );
  AOI21X2 U3293 ( .A0(mem_rdata[17]), .A1(n3900), .B0(n401), .Y(n227) );
  OAI22XL U3294 ( .A0(n3886), .A1(n4161), .B0(n3301), .B1(n3884), .Y(n401) );
  AOI21X2 U3295 ( .A0(mem_rdata[18]), .A1(n3900), .B0(n403), .Y(n228) );
  OAI22XL U3296 ( .A0(n3886), .A1(n4160), .B0(n3302), .B1(n3884), .Y(n403) );
  AOI21X2 U3297 ( .A0(mem_rdata[20]), .A1(n3899), .B0(n407), .Y(n230) );
  OAI22XL U3298 ( .A0(n3886), .A1(n4158), .B0(n3303), .B1(n3884), .Y(n407) );
  AOI21X2 U3299 ( .A0(mem_rdata[21]), .A1(n3899), .B0(n409), .Y(n231) );
  OAI22XL U3300 ( .A0(n3886), .A1(n4157), .B0(n3304), .B1(n3884), .Y(n409) );
  AOI21X2 U3301 ( .A0(mem_rdata[22]), .A1(n3899), .B0(n411), .Y(n232) );
  OAI22XL U3302 ( .A0(n3886), .A1(n4156), .B0(n3305), .B1(n3884), .Y(n411) );
  AOI21X2 U3303 ( .A0(mem_rdata[23]), .A1(n3899), .B0(n413), .Y(n233) );
  OAI22XL U3304 ( .A0(n3886), .A1(n4155), .B0(n3306), .B1(n3884), .Y(n413) );
  AOI21X2 U3305 ( .A0(mem_rdata[33]), .A1(n3898), .B0(n435), .Y(n243) );
  OAI22XL U3306 ( .A0(n4177), .A1(n3879), .B0(n3255), .B1(n3877), .Y(n435) );
  AOI21X2 U3307 ( .A0(mem_rdata[34]), .A1(n3898), .B0(n436), .Y(n244) );
  OAI22XL U3308 ( .A0(n4176), .A1(n3879), .B0(n3256), .B1(n3877), .Y(n436) );
  AOI21X2 U3309 ( .A0(mem_rdata[35]), .A1(n3898), .B0(n437), .Y(n245) );
  OAI22XL U3310 ( .A0(n4175), .A1(n3879), .B0(n3257), .B1(n3877), .Y(n437) );
  OAI22XL U3311 ( .A0(n4174), .A1(n3879), .B0(n3258), .B1(n3877), .Y(n438) );
  AOI21X2 U3312 ( .A0(mem_rdata[37]), .A1(n3898), .B0(n439), .Y(n247) );
  OAI22XL U3313 ( .A0(n4173), .A1(n3879), .B0(n3259), .B1(n3877), .Y(n439) );
  AOI21X2 U3314 ( .A0(mem_rdata[38]), .A1(n3898), .B0(n440), .Y(n248) );
  OAI22XL U3315 ( .A0(n4172), .A1(n3879), .B0(n3260), .B1(n3877), .Y(n440) );
  AOI21X2 U3316 ( .A0(mem_rdata[39]), .A1(n3898), .B0(n441), .Y(n249) );
  OAI22XL U3317 ( .A0(n4171), .A1(n3879), .B0(n3261), .B1(n3877), .Y(n441) );
  AOI21X2 U3318 ( .A0(mem_rdata[40]), .A1(n3898), .B0(n442), .Y(n250) );
  OAI22XL U3319 ( .A0(n4170), .A1(n3879), .B0(n3262), .B1(n3877), .Y(n442) );
  AOI21X2 U3320 ( .A0(mem_rdata[41]), .A1(n3898), .B0(n443), .Y(n251) );
  OAI22XL U3321 ( .A0(n4169), .A1(n3879), .B0(n3263), .B1(n3877), .Y(n443) );
  AOI21X2 U3322 ( .A0(mem_rdata[42]), .A1(n3898), .B0(n444), .Y(n252) );
  OAI22XL U3323 ( .A0(n4168), .A1(n3879), .B0(n3264), .B1(n3877), .Y(n444) );
  AOI21X2 U3324 ( .A0(mem_rdata[43]), .A1(n3897), .B0(n445), .Y(n253) );
  OAI22XL U3325 ( .A0(n4167), .A1(n3879), .B0(n3265), .B1(n3877), .Y(n445) );
  AOI21X2 U3326 ( .A0(mem_rdata[44]), .A1(n3897), .B0(n446), .Y(n254) );
  AOI21X2 U3327 ( .A0(mem_rdata[45]), .A1(n3897), .B0(n447), .Y(n255) );
  OAI22XL U3328 ( .A0(n4165), .A1(n3880), .B0(n3267), .B1(n3878), .Y(n447) );
  AOI21X2 U3329 ( .A0(mem_rdata[46]), .A1(n3897), .B0(n448), .Y(n256) );
  OAI22XL U3330 ( .A0(n4164), .A1(n3880), .B0(n3268), .B1(n3878), .Y(n448) );
  AOI21X2 U3331 ( .A0(mem_rdata[47]), .A1(n3897), .B0(n449), .Y(n257) );
  OAI22XL U3332 ( .A0(n4163), .A1(n3880), .B0(n3269), .B1(n3878), .Y(n449) );
  AOI21X2 U3333 ( .A0(mem_rdata[48]), .A1(n3897), .B0(n450), .Y(n258) );
  OAI22XL U3334 ( .A0(n4162), .A1(n3880), .B0(n3270), .B1(n3878), .Y(n450) );
  AOI21X2 U3335 ( .A0(mem_rdata[49]), .A1(n3897), .B0(n451), .Y(n259) );
  OAI22XL U3336 ( .A0(n4161), .A1(n3880), .B0(n3271), .B1(n3878), .Y(n451) );
  AOI21X2 U3337 ( .A0(mem_rdata[50]), .A1(n3897), .B0(n452), .Y(n260) );
  OAI22XL U3338 ( .A0(n4160), .A1(n3880), .B0(n3272), .B1(n3878), .Y(n452) );
  AOI21X2 U3339 ( .A0(mem_rdata[51]), .A1(n3897), .B0(n453), .Y(n261) );
  OAI22XL U3340 ( .A0(n4159), .A1(n3880), .B0(n3273), .B1(n3878), .Y(n453) );
  AOI21X2 U3341 ( .A0(mem_rdata[52]), .A1(n3897), .B0(n454), .Y(n262) );
  OAI22XL U3342 ( .A0(n4158), .A1(n3880), .B0(n3274), .B1(n3878), .Y(n454) );
  AOI21X2 U3343 ( .A0(mem_rdata[53]), .A1(n3897), .B0(n455), .Y(n263) );
  OAI22XL U3344 ( .A0(n4157), .A1(n3880), .B0(n3275), .B1(n3878), .Y(n455) );
  AOI21X2 U3345 ( .A0(mem_rdata[54]), .A1(n3893), .B0(n456), .Y(n264) );
  OAI22XL U3346 ( .A0(n4156), .A1(n3880), .B0(n3276), .B1(n3878), .Y(n456) );
  AOI21X2 U3347 ( .A0(mem_rdata[55]), .A1(n3893), .B0(n457), .Y(n265) );
  OAI22XL U3348 ( .A0(n4155), .A1(n3880), .B0(n3277), .B1(n3878), .Y(n457) );
  AOI21X2 U3349 ( .A0(mem_rdata[64]), .A1(n3893), .B0(n466), .Y(n274) );
  OAI22XL U3350 ( .A0(n4178), .A1(n3874), .B0(n3192), .B1(n3087), .Y(n466) );
  AOI21X2 U3351 ( .A0(mem_rdata[65]), .A1(n3893), .B0(n469), .Y(n275) );
  OAI22XL U3352 ( .A0(n4177), .A1(n3874), .B0(n3193), .B1(n3087), .Y(n469) );
  AOI21X2 U3353 ( .A0(mem_rdata[66]), .A1(n3899), .B0(n470), .Y(n276) );
  OAI22XL U3354 ( .A0(n4176), .A1(n3874), .B0(n3194), .B1(n3087), .Y(n470) );
  AOI21X2 U3355 ( .A0(mem_rdata[67]), .A1(n3898), .B0(n471), .Y(n277) );
  OAI22XL U3356 ( .A0(n4175), .A1(n3874), .B0(n3195), .B1(n3087), .Y(n471) );
  AOI21X2 U3357 ( .A0(mem_rdata[68]), .A1(n3897), .B0(n472), .Y(n278) );
  OAI22XL U3358 ( .A0(n4174), .A1(n3874), .B0(n3196), .B1(n3087), .Y(n472) );
  AOI21X2 U3359 ( .A0(mem_rdata[69]), .A1(n3893), .B0(n473), .Y(n279) );
  OAI22XL U3360 ( .A0(n4173), .A1(n3874), .B0(n3197), .B1(n3087), .Y(n473) );
  AOI21X2 U3361 ( .A0(mem_rdata[70]), .A1(n3901), .B0(n474), .Y(n280) );
  OAI22XL U3362 ( .A0(n4172), .A1(n3874), .B0(n3198), .B1(n3087), .Y(n474) );
  AOI21X2 U3363 ( .A0(mem_rdata[71]), .A1(n3893), .B0(n475), .Y(n281) );
  OAI22XL U3364 ( .A0(n4171), .A1(n3874), .B0(n3206), .B1(n3087), .Y(n475) );
  AOI21X2 U3365 ( .A0(mem_rdata[72]), .A1(n3902), .B0(n476), .Y(n282) );
  OAI22XL U3366 ( .A0(n4170), .A1(n3874), .B0(n3207), .B1(n3087), .Y(n476) );
  AOI21X2 U3367 ( .A0(mem_rdata[73]), .A1(n3900), .B0(n477), .Y(n283) );
  OAI22XL U3368 ( .A0(n4169), .A1(n3874), .B0(n3208), .B1(n3087), .Y(n477) );
  AOI21X2 U3369 ( .A0(mem_rdata[74]), .A1(n3899), .B0(n478), .Y(n284) );
  OAI22XL U3370 ( .A0(n4168), .A1(n3874), .B0(n3209), .B1(n3087), .Y(n478) );
  AOI21X2 U3371 ( .A0(mem_rdata[75]), .A1(n3898), .B0(n479), .Y(n285) );
  OAI22XL U3372 ( .A0(n4167), .A1(n3874), .B0(n3210), .B1(n3087), .Y(n479) );
  AOI21X2 U3373 ( .A0(mem_rdata[76]), .A1(n3893), .B0(n480), .Y(n286) );
  OAI22XL U3374 ( .A0(n4166), .A1(n3875), .B0(n3211), .B1(n3087), .Y(n480) );
  AOI21X2 U3375 ( .A0(mem_rdata[77]), .A1(n351), .B0(n481), .Y(n287) );
  OAI22XL U3376 ( .A0(n4165), .A1(n3875), .B0(n3212), .B1(n3087), .Y(n481) );
  AOI21X2 U3377 ( .A0(mem_rdata[78]), .A1(n3894), .B0(n482), .Y(n288) );
  OAI22XL U3378 ( .A0(n4164), .A1(n3875), .B0(n3213), .B1(n3087), .Y(n482) );
  AOI21X2 U3379 ( .A0(mem_rdata[79]), .A1(n3896), .B0(n483), .Y(n289) );
  OAI22XL U3380 ( .A0(n4163), .A1(n3875), .B0(n3214), .B1(n3087), .Y(n483) );
  AOI21X2 U3381 ( .A0(mem_rdata[80]), .A1(n3899), .B0(n484), .Y(n290) );
  OAI22XL U3382 ( .A0(n4162), .A1(n3875), .B0(n3215), .B1(n3087), .Y(n484) );
  AOI21X2 U3383 ( .A0(mem_rdata[81]), .A1(n3897), .B0(n485), .Y(n291) );
  OAI22XL U3384 ( .A0(n4161), .A1(n3875), .B0(n3216), .B1(n3087), .Y(n485) );
  AOI21X2 U3385 ( .A0(mem_rdata[82]), .A1(n3901), .B0(n486), .Y(n292) );
  OAI22XL U3386 ( .A0(n4160), .A1(n3875), .B0(n3217), .B1(n3087), .Y(n486) );
  AOI21X2 U3387 ( .A0(mem_rdata[83]), .A1(n3902), .B0(n487), .Y(n293) );
  OAI22XL U3388 ( .A0(n4159), .A1(n3875), .B0(n3218), .B1(n3087), .Y(n487) );
  AOI21X2 U3389 ( .A0(mem_rdata[84]), .A1(n3900), .B0(n488), .Y(n294) );
  OAI22XL U3390 ( .A0(n4158), .A1(n3875), .B0(n3219), .B1(n3087), .Y(n488) );
  AOI21X2 U3391 ( .A0(mem_rdata[85]), .A1(n3895), .B0(n489), .Y(n295) );
  OAI22XL U3392 ( .A0(n4157), .A1(n3875), .B0(n3220), .B1(n3087), .Y(n489) );
  AOI21X2 U3393 ( .A0(mem_rdata[86]), .A1(n3894), .B0(n490), .Y(n296) );
  OAI22XL U3394 ( .A0(n4156), .A1(n3875), .B0(n3221), .B1(n3087), .Y(n490) );
  AOI21X2 U3395 ( .A0(mem_rdata[87]), .A1(n3896), .B0(n491), .Y(n297) );
  OAI22XL U3396 ( .A0(n4155), .A1(n3875), .B0(n3222), .B1(n3087), .Y(n491) );
  AOI21X2 U3397 ( .A0(mem_rdata[96]), .A1(n3896), .B0(n500), .Y(n306) );
  OAI22XL U3398 ( .A0(n3890), .A1(n4178), .B0(n3278), .B1(n3075), .Y(n500) );
  AOI21X2 U3399 ( .A0(mem_rdata[97]), .A1(n3896), .B0(n501), .Y(n307) );
  OAI22XL U3400 ( .A0(n3890), .A1(n4177), .B0(n3279), .B1(n3075), .Y(n501) );
  AOI21X2 U3401 ( .A0(mem_rdata[98]), .A1(n3896), .B0(n502), .Y(n308) );
  OAI22XL U3402 ( .A0(n3890), .A1(n4176), .B0(n3280), .B1(n3075), .Y(n502) );
  AOI21X2 U3403 ( .A0(mem_rdata[99]), .A1(n3896), .B0(n503), .Y(n309) );
  OAI22XL U3404 ( .A0(n3890), .A1(n4175), .B0(n3281), .B1(n3075), .Y(n503) );
  AOI21X2 U3405 ( .A0(mem_rdata[100]), .A1(n3896), .B0(n504), .Y(n310) );
  OAI22XL U3406 ( .A0(n3890), .A1(n4174), .B0(n3282), .B1(n3075), .Y(n504) );
  AOI21X2 U3407 ( .A0(mem_rdata[101]), .A1(n3896), .B0(n505), .Y(n311) );
  OAI22XL U3408 ( .A0(n3890), .A1(n4173), .B0(n3283), .B1(n3075), .Y(n505) );
  AOI21X2 U3409 ( .A0(mem_rdata[102]), .A1(n3895), .B0(n506), .Y(n312) );
  OAI22XL U3410 ( .A0(n3890), .A1(n4172), .B0(n3284), .B1(n3075), .Y(n506) );
  AOI21X2 U3411 ( .A0(mem_rdata[103]), .A1(n3895), .B0(n507), .Y(n313) );
  OAI22XL U3412 ( .A0(n3890), .A1(n4171), .B0(n3285), .B1(n3075), .Y(n507) );
  AOI21X2 U3413 ( .A0(mem_rdata[104]), .A1(n3895), .B0(n508), .Y(n314) );
  OAI22XL U3414 ( .A0(n3890), .A1(n4170), .B0(n3286), .B1(n3075), .Y(n508) );
  AOI21X2 U3415 ( .A0(mem_rdata[105]), .A1(n3895), .B0(n509), .Y(n315) );
  OAI22XL U3416 ( .A0(n3890), .A1(n4169), .B0(n3287), .B1(n3075), .Y(n509) );
  AOI21X2 U3417 ( .A0(mem_rdata[106]), .A1(n3895), .B0(n510), .Y(n316) );
  OAI22XL U3418 ( .A0(n3891), .A1(n4168), .B0(n3288), .B1(n3075), .Y(n510) );
  AOI21X2 U3419 ( .A0(mem_rdata[107]), .A1(n3895), .B0(n511), .Y(n317) );
  OAI22XL U3420 ( .A0(n3891), .A1(n4167), .B0(n3224), .B1(n3075), .Y(n511) );
  AOI21X2 U3421 ( .A0(mem_rdata[108]), .A1(n3895), .B0(n512), .Y(n318) );
  OAI22XL U3422 ( .A0(n3891), .A1(n4166), .B0(n3225), .B1(n3075), .Y(n512) );
  AOI21X2 U3423 ( .A0(mem_rdata[109]), .A1(n3895), .B0(n513), .Y(n319) );
  OAI22XL U3424 ( .A0(n3891), .A1(n4165), .B0(n3226), .B1(n3075), .Y(n513) );
  AOI21X2 U3425 ( .A0(mem_rdata[110]), .A1(n3895), .B0(n514), .Y(n320) );
  OAI22XL U3426 ( .A0(n3891), .A1(n4164), .B0(n3227), .B1(n3075), .Y(n514) );
  AOI21X2 U3427 ( .A0(mem_rdata[111]), .A1(n3895), .B0(n515), .Y(n321) );
  OAI22XL U3428 ( .A0(n3891), .A1(n4163), .B0(n3228), .B1(n3075), .Y(n515) );
  AOI21X2 U3429 ( .A0(mem_rdata[112]), .A1(n3895), .B0(n516), .Y(n322) );
  OAI22XL U3430 ( .A0(n3891), .A1(n4162), .B0(n3229), .B1(n3075), .Y(n516) );
  AOI21X2 U3431 ( .A0(mem_rdata[113]), .A1(n3895), .B0(n517), .Y(n323) );
  OAI22XL U3432 ( .A0(n3891), .A1(n4161), .B0(n3230), .B1(n3075), .Y(n517) );
  AOI21X2 U3433 ( .A0(mem_rdata[114]), .A1(n3894), .B0(n518), .Y(n324) );
  OAI22XL U3434 ( .A0(n3891), .A1(n4160), .B0(n3231), .B1(n3075), .Y(n518) );
  AOI21X2 U3435 ( .A0(mem_rdata[115]), .A1(n3894), .B0(n519), .Y(n325) );
  OAI22XL U3436 ( .A0(n3891), .A1(n4159), .B0(n3232), .B1(n3075), .Y(n519) );
  AOI21X2 U3437 ( .A0(mem_rdata[116]), .A1(n3894), .B0(n520), .Y(n326) );
  OAI22XL U3438 ( .A0(n3891), .A1(n4158), .B0(n3233), .B1(n3075), .Y(n520) );
  AOI21X2 U3439 ( .A0(mem_rdata[117]), .A1(n3894), .B0(n521), .Y(n327) );
  OAI22XL U3440 ( .A0(n3891), .A1(n4157), .B0(n3234), .B1(n3075), .Y(n521) );
  AOI21X2 U3441 ( .A0(mem_rdata[126]), .A1(n3894), .B0(n352), .Y(n178) );
  OAI22XL U3442 ( .A0(n3890), .A1(n4148), .B0(n3375), .B1(n3075), .Y(n352) );
  OAI22XL U3443 ( .A0(n572), .A1(n3931), .B0(n3080), .B1(n3953), .Y(n1812) );
  OAI22XL U3444 ( .A0(n573), .A1(n3931), .B0(n211), .B1(n3944), .Y(n1813) );
  OAI22XL U3445 ( .A0(n574), .A1(n3931), .B0(n3081), .B1(n3956), .Y(n1814) );
  OAI22XL U3446 ( .A0(n575), .A1(n3931), .B0(n3079), .B1(n3947), .Y(n1815) );
  OAI22XL U3447 ( .A0(n576), .A1(n3931), .B0(n3078), .B1(n3945), .Y(n1816) );
  OAI22XL U3448 ( .A0(n577), .A1(n3931), .B0(n3077), .B1(n3945), .Y(n1817) );
  OAI22XL U3449 ( .A0(n578), .A1(n3931), .B0(n3076), .B1(n3945), .Y(n1818) );
  OAI22XL U3450 ( .A0(n579), .A1(n3931), .B0(n3086), .B1(n3945), .Y(n1819) );
  OAI22XL U3451 ( .A0(n580), .A1(n3931), .B0(n3085), .B1(n3945), .Y(n1820) );
  OAI22XL U3452 ( .A0(n581), .A1(n3931), .B0(n3084), .B1(n3945), .Y(n1821) );
  OAI22XL U3453 ( .A0(n582), .A1(n3931), .B0(n3083), .B1(n3945), .Y(n1822) );
  OAI22XL U3454 ( .A0(n583), .A1(n3931), .B0(n3082), .B1(n3945), .Y(n1823) );
  OAI22XL U3455 ( .A0(n584), .A1(n3932), .B0(n222), .B1(n3946), .Y(n1824) );
  OAI22XL U3456 ( .A0(n585), .A1(n3932), .B0(n223), .B1(n3946), .Y(n1825) );
  OAI22XL U3457 ( .A0(n586), .A1(n3932), .B0(n3130), .B1(n3946), .Y(n1826) );
  OAI22XL U3458 ( .A0(n587), .A1(n3932), .B0(n3129), .B1(n3946), .Y(n1827) );
  OAI22XL U3459 ( .A0(n588), .A1(n3932), .B0(n3128), .B1(n3946), .Y(n1828) );
  OAI22XL U3460 ( .A0(n589), .A1(n3932), .B0(n3127), .B1(n3946), .Y(n1829) );
  OAI22XL U3461 ( .A0(n590), .A1(n3932), .B0(n3126), .B1(n3946), .Y(n1830) );
  OAI22XL U3462 ( .A0(n591), .A1(n3932), .B0(n229), .B1(n3946), .Y(n1831) );
  OAI22XL U3463 ( .A0(n592), .A1(n3932), .B0(n3134), .B1(n3946), .Y(n1832) );
  OAI22XL U3464 ( .A0(n593), .A1(n3932), .B0(n3133), .B1(n3946), .Y(n1833) );
  OAI22XL U3465 ( .A0(n594), .A1(n3932), .B0(n3132), .B1(n3946), .Y(n1834) );
  OAI22XL U3466 ( .A0(n595), .A1(n3932), .B0(n3131), .B1(n3954), .Y(n1835) );
  OAI22XL U3467 ( .A0(n596), .A1(n3933), .B0(n3073), .B1(n3956), .Y(n1836) );
  OAI22XL U3468 ( .A0(n597), .A1(n3933), .B0(n3067), .B1(n3953), .Y(n1837) );
  OAI22XL U3469 ( .A0(n598), .A1(n3933), .B0(n3064), .B1(n3954), .Y(n1838) );
  OAI22XL U3470 ( .A0(n599), .A1(n3933), .B0(n3070), .B1(n3956), .Y(n1839) );
  OAI22XL U3471 ( .A0(n600), .A1(n3933), .B0(n3061), .B1(n3953), .Y(n1840) );
  OAI22XL U3472 ( .A0(n601), .A1(n3933), .B0(n3058), .B1(n3954), .Y(n1841) );
  OAI22XL U3473 ( .A0(n602), .A1(n3933), .B0(n3055), .B1(n3956), .Y(n1842) );
  OAI22XL U3474 ( .A0(n603), .A1(n3933), .B0(n3053), .B1(n3953), .Y(n1843) );
  OAI22XL U3475 ( .A0(n605), .A1(n3933), .B0(n3125), .B1(n3954), .Y(n1845) );
  OAI22XL U3476 ( .A0(n606), .A1(n3933), .B0(n3124), .B1(n3947), .Y(n1846) );
  OAI22XL U3477 ( .A0(n607), .A1(n3933), .B0(n3123), .B1(n3947), .Y(n1847) );
  OAI22XL U3478 ( .A0(n609), .A1(n3934), .B0(n3122), .B1(n3947), .Y(n1849) );
  OAI22XL U3479 ( .A0(n610), .A1(n3934), .B0(n3121), .B1(n3947), .Y(n1850) );
  OAI22XL U3480 ( .A0(n611), .A1(n3934), .B0(n3120), .B1(n3947), .Y(n1851) );
  OAI22XL U3481 ( .A0(n612), .A1(n3934), .B0(n3119), .B1(n3947), .Y(n1852) );
  OAI22XL U3482 ( .A0(n613), .A1(n3934), .B0(n3118), .B1(n3947), .Y(n1853) );
  OAI22XL U3483 ( .A0(n614), .A1(n3934), .B0(n3117), .B1(n3947), .Y(n1854) );
  OAI22XL U3484 ( .A0(n615), .A1(n3934), .B0(n3116), .B1(n3947), .Y(n1855) );
  OAI22XL U3485 ( .A0(n616), .A1(n3934), .B0(n3115), .B1(n3947), .Y(n1856) );
  OAI22XL U3486 ( .A0(n617), .A1(n3934), .B0(n3114), .B1(n3948), .Y(n1857) );
  OAI22XL U3487 ( .A0(n618), .A1(n3934), .B0(n3113), .B1(n3948), .Y(n1858) );
  OAI22XL U3488 ( .A0(n619), .A1(n3934), .B0(n3112), .B1(n3948), .Y(n1859) );
  OAI22XL U3489 ( .A0(n620), .A1(n3935), .B0(n3111), .B1(n3948), .Y(n1860) );
  OAI22XL U3490 ( .A0(n621), .A1(n3935), .B0(n3110), .B1(n3948), .Y(n1861) );
  OAI22XL U3491 ( .A0(n622), .A1(n3935), .B0(n3109), .B1(n3948), .Y(n1862) );
  OAI22XL U3492 ( .A0(n623), .A1(n3935), .B0(n3108), .B1(n3948), .Y(n1863) );
  OAI22XL U3493 ( .A0(n624), .A1(n3935), .B0(n3107), .B1(n3948), .Y(n1864) );
  OAI22XL U3494 ( .A0(n625), .A1(n3935), .B0(n3106), .B1(n3948), .Y(n1865) );
  OAI22XL U3495 ( .A0(n626), .A1(n3935), .B0(n3105), .B1(n3948), .Y(n1866) );
  OAI22XL U3496 ( .A0(n627), .A1(n3935), .B0(n3104), .B1(n3948), .Y(n1867) );
  OAI22XL U3497 ( .A0(n628), .A1(n3935), .B0(n3103), .B1(n3949), .Y(n1868) );
  OAI22XL U3498 ( .A0(n629), .A1(n3935), .B0(n3102), .B1(n3949), .Y(n1869) );
  OAI22XL U3499 ( .A0(n630), .A1(n3935), .B0(n3089), .B1(n3949), .Y(n1870) );
  OAI22XL U3500 ( .A0(n631), .A1(n3935), .B0(n3101), .B1(n3949), .Y(n1871) );
  OAI22XL U3501 ( .A0(n632), .A1(n3936), .B0(n3100), .B1(n3949), .Y(n1872) );
  OAI22XL U3502 ( .A0(n633), .A1(n3936), .B0(n3099), .B1(n3949), .Y(n1873) );
  OAI22XL U3503 ( .A0(n634), .A1(n3936), .B0(n3098), .B1(n3949), .Y(n1874) );
  OAI22XL U3504 ( .A0(n635), .A1(n3936), .B0(n3088), .B1(n3949), .Y(n1875) );
  OAI22XL U3505 ( .A0(n636), .A1(n3936), .B0(n3152), .B1(n3949), .Y(n1876) );
  OAI22XL U3506 ( .A0(n637), .A1(n3936), .B0(n3151), .B1(n3949), .Y(n1877) );
  OAI22XL U3507 ( .A0(n638), .A1(n3936), .B0(n3168), .B1(n3949), .Y(n1878) );
  OAI22XL U3508 ( .A0(n639), .A1(n3936), .B0(n3170), .B1(n3950), .Y(n1879) );
  OAI22XL U3509 ( .A0(n640), .A1(n3936), .B0(n3159), .B1(n3950), .Y(n1880) );
  OAI22XL U3510 ( .A0(n641), .A1(n3936), .B0(n3150), .B1(n3950), .Y(n1881) );
  OAI22XL U3511 ( .A0(n642), .A1(n3936), .B0(n3161), .B1(n3950), .Y(n1882) );
  OAI22XL U3512 ( .A0(n643), .A1(n3936), .B0(n3149), .B1(n3950), .Y(n1883) );
  OAI22XL U3513 ( .A0(n644), .A1(n3937), .B0(n3163), .B1(n3950), .Y(n1884) );
  OAI22XL U3514 ( .A0(n645), .A1(n3937), .B0(n3165), .B1(n3950), .Y(n1885) );
  OAI22XL U3515 ( .A0(n646), .A1(n3937), .B0(n3167), .B1(n3950), .Y(n1886) );
  OAI22XL U3516 ( .A0(n647), .A1(n3937), .B0(n3169), .B1(n3950), .Y(n1887) );
  OAI22XL U3517 ( .A0(n648), .A1(n3937), .B0(n3148), .B1(n3950), .Y(n1888) );
  OAI22XL U3518 ( .A0(n649), .A1(n3937), .B0(n3147), .B1(n3950), .Y(n1889) );
  OAI22XL U3519 ( .A0(n650), .A1(n3937), .B0(n3158), .B1(n3951), .Y(n1890) );
  OAI22XL U3520 ( .A0(n651), .A1(n3937), .B0(n3157), .B1(n3951), .Y(n1891) );
  OAI22XL U3521 ( .A0(n652), .A1(n3937), .B0(n3166), .B1(n3951), .Y(n1892) );
  OAI22XL U3522 ( .A0(n653), .A1(n3937), .B0(n3156), .B1(n3951), .Y(n1893) );
  OAI22XL U3523 ( .A0(n654), .A1(n3937), .B0(n3160), .B1(n3951), .Y(n1894) );
  OAI22XL U3524 ( .A0(n655), .A1(n3937), .B0(n3162), .B1(n3951), .Y(n1895) );
  OAI22XL U3525 ( .A0(n656), .A1(n3938), .B0(n3164), .B1(n3951), .Y(n1896) );
  OAI22XL U3526 ( .A0(n657), .A1(n3938), .B0(n3155), .B1(n3951), .Y(n1897) );
  OAI22XL U3527 ( .A0(n658), .A1(n3938), .B0(n3154), .B1(n3951), .Y(n1898) );
  OAI22XL U3528 ( .A0(n659), .A1(n3938), .B0(n3153), .B1(n3951), .Y(n1899) );
  OAI22XL U3529 ( .A0(n660), .A1(n3938), .B0(n3097), .B1(n3951), .Y(n1900) );
  OAI22XL U3530 ( .A0(n661), .A1(n3938), .B0(n3093), .B1(n3952), .Y(n1901) );
  OAI22XL U3531 ( .A0(n662), .A1(n3938), .B0(n3092), .B1(n3952), .Y(n1902) );
  OAI22XL U3532 ( .A0(n663), .A1(n3938), .B0(n3091), .B1(n3952), .Y(n1903) );
  OAI22XL U3533 ( .A0(n664), .A1(n3938), .B0(n3090), .B1(n3952), .Y(n1904) );
  OAI22XL U3534 ( .A0(n665), .A1(n3938), .B0(n3096), .B1(n3952), .Y(n1905) );
  OAI22XL U3535 ( .A0(n666), .A1(n3938), .B0(n3095), .B1(n3952), .Y(n1906) );
  OAI22XL U3536 ( .A0(n667), .A1(n3938), .B0(n3094), .B1(n3952), .Y(n1907) );
  OAI22XL U3537 ( .A0(n668), .A1(n3939), .B0(n3179), .B1(n3952), .Y(n1908) );
  OAI22XL U3538 ( .A0(n669), .A1(n3939), .B0(n3178), .B1(n3952), .Y(n1909) );
  OAI22XL U3539 ( .A0(n670), .A1(n3939), .B0(n3177), .B1(n3952), .Y(n1910) );
  OAI22XL U3540 ( .A0(n671), .A1(n3939), .B0(n3176), .B1(n3952), .Y(n1911) );
  OAI22XL U3541 ( .A0(n672), .A1(n3939), .B0(n3187), .B1(n3953), .Y(n1912) );
  OAI22XL U3542 ( .A0(n673), .A1(n3939), .B0(n3186), .B1(n3953), .Y(n1913) );
  OAI22XL U3543 ( .A0(n674), .A1(n3939), .B0(n3185), .B1(n3953), .Y(n1914) );
  OAI22XL U3544 ( .A0(n675), .A1(n3939), .B0(n3184), .B1(n3953), .Y(n1915) );
  OAI22XL U3545 ( .A0(n676), .A1(n3939), .B0(n3183), .B1(n3953), .Y(n1916) );
  OAI22XL U3546 ( .A0(n677), .A1(n3939), .B0(n3182), .B1(n3953), .Y(n1917) );
  OAI22XL U3547 ( .A0(n678), .A1(n3939), .B0(n3146), .B1(n3953), .Y(n1918) );
  OAI22XL U3548 ( .A0(n679), .A1(n3939), .B0(n3145), .B1(n3953), .Y(n1919) );
  OAI22XL U3549 ( .A0(n680), .A1(n3940), .B0(n3144), .B1(n3953), .Y(n1920) );
  OAI22XL U3550 ( .A0(n681), .A1(n3940), .B0(n3143), .B1(n3953), .Y(n1921) );
  OAI22XL U3551 ( .A0(n682), .A1(n3940), .B0(n3142), .B1(n3953), .Y(n1922) );
  OAI22XL U3552 ( .A0(n683), .A1(n3940), .B0(n3139), .B1(n3950), .Y(n1923) );
  OAI22XL U3553 ( .A0(n684), .A1(n3940), .B0(n3138), .B1(n3951), .Y(n1924) );
  OAI22XL U3554 ( .A0(n685), .A1(n3940), .B0(n3137), .B1(n3949), .Y(n1925) );
  OAI22XL U3555 ( .A0(n686), .A1(n3940), .B0(n3136), .B1(n3948), .Y(n1926) );
  OAI22XL U3556 ( .A0(n687), .A1(n3940), .B0(n3141), .B1(n3950), .Y(n1927) );
  OAI22XL U3557 ( .A0(n688), .A1(n3940), .B0(n3135), .B1(n3951), .Y(n1928) );
  OAI22XL U3558 ( .A0(n689), .A1(n3940), .B0(n3140), .B1(n3949), .Y(n1929) );
  OAI22XL U3559 ( .A0(n690), .A1(n3940), .B0(n3172), .B1(n3948), .Y(n1930) );
  OAI22XL U3560 ( .A0(n691), .A1(n3940), .B0(n3180), .B1(n3950), .Y(n1931) );
  OAI22XL U3561 ( .A0(n692), .A1(n3941), .B0(n3173), .B1(n3951), .Y(n1932) );
  OAI22XL U3562 ( .A0(n693), .A1(n3941), .B0(n3171), .B1(n3949), .Y(n1933) );
  OAI22XL U3563 ( .A0(n694), .A1(n3941), .B0(n3189), .B1(n3954), .Y(n1934) );
  OAI22XL U3564 ( .A0(n695), .A1(n3941), .B0(n3188), .B1(n3954), .Y(n1935) );
  OAI22XL U3565 ( .A0(n696), .A1(n3941), .B0(n3175), .B1(n3954), .Y(n1936) );
  OAI22XL U3566 ( .A0(n697), .A1(n3941), .B0(n3181), .B1(n3954), .Y(n1937) );
  OAI22XL U3567 ( .A0(n698), .A1(n3941), .B0(n3174), .B1(n3954), .Y(n1938) );
  OAI22XL U3568 ( .A0(n727), .A1(n3903), .B0(n3080), .B1(n3928), .Y(n1967) );
  OAI22XL U3569 ( .A0(n728), .A1(n3903), .B0(n211), .B1(n3926), .Y(n1968) );
  OAI22XL U3570 ( .A0(n729), .A1(n3903), .B0(n3081), .B1(n3917), .Y(n1969) );
  OAI22XL U3571 ( .A0(n730), .A1(n3903), .B0(n3079), .B1(n3927), .Y(n1970) );
  OAI22XL U3572 ( .A0(n731), .A1(n3903), .B0(n3078), .B1(n3916), .Y(n1971) );
  OAI22XL U3573 ( .A0(n732), .A1(n3903), .B0(n3077), .B1(n3916), .Y(n1972) );
  OAI22XL U3574 ( .A0(n733), .A1(n3903), .B0(n3076), .B1(n3916), .Y(n1973) );
  OAI22XL U3575 ( .A0(n734), .A1(n3903), .B0(n3086), .B1(n3916), .Y(n1974) );
  OAI22XL U3576 ( .A0(n735), .A1(n3903), .B0(n3085), .B1(n3916), .Y(n1975) );
  OAI22XL U3577 ( .A0(n736), .A1(n3903), .B0(n3084), .B1(n3916), .Y(n1976) );
  OAI22XL U3578 ( .A0(n737), .A1(n3903), .B0(n3083), .B1(n3916), .Y(n1977) );
  OAI22XL U3579 ( .A0(n738), .A1(n3903), .B0(n3082), .B1(n3916), .Y(n1978) );
  OAI22XL U3580 ( .A0(n739), .A1(n3904), .B0(n222), .B1(n3917), .Y(n1979) );
  OAI22XL U3581 ( .A0(n740), .A1(n3904), .B0(n223), .B1(n3917), .Y(n1980) );
  OAI22XL U3582 ( .A0(n741), .A1(n3904), .B0(n3130), .B1(n3917), .Y(n1981) );
  OAI22XL U3583 ( .A0(n742), .A1(n3904), .B0(n3129), .B1(n3917), .Y(n1982) );
  OAI22XL U3584 ( .A0(n743), .A1(n3904), .B0(n3128), .B1(n3917), .Y(n1983) );
  OAI22XL U3585 ( .A0(n744), .A1(n3904), .B0(n3127), .B1(n3917), .Y(n1984) );
  OAI22XL U3586 ( .A0(n745), .A1(n3904), .B0(n3126), .B1(n3917), .Y(n1985) );
  OAI22XL U3587 ( .A0(n746), .A1(n3904), .B0(n229), .B1(n3917), .Y(n1986) );
  OAI22XL U3588 ( .A0(n747), .A1(n3904), .B0(n3134), .B1(n3917), .Y(n1987) );
  OAI22XL U3589 ( .A0(n748), .A1(n3904), .B0(n3133), .B1(n3917), .Y(n1988) );
  OAI22XL U3590 ( .A0(n749), .A1(n3904), .B0(n3132), .B1(n3917), .Y(n1989) );
  OAI22XL U3591 ( .A0(n750), .A1(n3904), .B0(n3131), .B1(n3918), .Y(n1990) );
  OAI22XL U3592 ( .A0(n751), .A1(n3905), .B0(n3074), .B1(n3918), .Y(n1991) );
  OAI22XL U3593 ( .A0(n752), .A1(n3905), .B0(n3068), .B1(n3918), .Y(n1992) );
  OAI22XL U3594 ( .A0(n753), .A1(n3905), .B0(n3065), .B1(n3918), .Y(n1993) );
  OAI22XL U3595 ( .A0(n754), .A1(n3905), .B0(n3070), .B1(n3918), .Y(n1994) );
  OAI22XL U3596 ( .A0(n755), .A1(n3905), .B0(n3061), .B1(n3918), .Y(n1995) );
  OAI22XL U3597 ( .A0(n756), .A1(n3905), .B0(n3058), .B1(n3918), .Y(n1996) );
  OAI22XL U3598 ( .A0(n757), .A1(n3905), .B0(n3055), .B1(n3918), .Y(n1997) );
  OAI22XL U3599 ( .A0(n758), .A1(n3905), .B0(n3053), .B1(n3918), .Y(n1998) );
  OAI22XL U3600 ( .A0(n759), .A1(n3905), .B0(n242), .B1(n3918), .Y(n1999) );
  OAI22XL U3601 ( .A0(n760), .A1(n3905), .B0(n3125), .B1(n3918), .Y(n2000) );
  OAI22XL U3602 ( .A0(n761), .A1(n3905), .B0(n3124), .B1(n3919), .Y(n2001) );
  OAI22XL U3603 ( .A0(n762), .A1(n3905), .B0(n3123), .B1(n3919), .Y(n2002) );
  OAI22XL U3604 ( .A0(n763), .A1(n3906), .B0(n246), .B1(n3919), .Y(n2003) );
  OAI22XL U3605 ( .A0(n764), .A1(n3906), .B0(n3122), .B1(n3919), .Y(n2004) );
  OAI22XL U3606 ( .A0(n765), .A1(n3906), .B0(n3121), .B1(n3919), .Y(n2005) );
  OAI22XL U3607 ( .A0(n766), .A1(n3906), .B0(n3120), .B1(n3919), .Y(n2006) );
  OAI22XL U3608 ( .A0(n767), .A1(n3906), .B0(n3119), .B1(n3919), .Y(n2007) );
  OAI22XL U3609 ( .A0(n768), .A1(n3906), .B0(n3118), .B1(n3919), .Y(n2008) );
  OAI22XL U3610 ( .A0(n769), .A1(n3906), .B0(n3117), .B1(n3919), .Y(n2009) );
  OAI22XL U3611 ( .A0(n770), .A1(n3906), .B0(n3116), .B1(n3919), .Y(n2010) );
  OAI22XL U3612 ( .A0(n771), .A1(n3906), .B0(n3115), .B1(n3919), .Y(n2011) );
  OAI22XL U3613 ( .A0(n772), .A1(n3906), .B0(n3114), .B1(n3920), .Y(n2012) );
  OAI22XL U3614 ( .A0(n773), .A1(n3906), .B0(n3113), .B1(n3920), .Y(n2013) );
  OAI22XL U3615 ( .A0(n774), .A1(n3906), .B0(n3112), .B1(n3920), .Y(n2014) );
  OAI22XL U3616 ( .A0(n775), .A1(n3907), .B0(n3111), .B1(n3920), .Y(n2015) );
  OAI22XL U3617 ( .A0(n776), .A1(n3907), .B0(n3110), .B1(n3920), .Y(n2016) );
  OAI22XL U3618 ( .A0(n777), .A1(n3907), .B0(n3109), .B1(n3920), .Y(n2017) );
  OAI22XL U3619 ( .A0(n778), .A1(n3907), .B0(n3108), .B1(n3920), .Y(n2018) );
  OAI22XL U3620 ( .A0(n779), .A1(n3907), .B0(n3107), .B1(n3920), .Y(n2019) );
  OAI22XL U3621 ( .A0(n780), .A1(n3907), .B0(n3106), .B1(n3920), .Y(n2020) );
  OAI22XL U3622 ( .A0(n781), .A1(n3907), .B0(n3105), .B1(n3920), .Y(n2021) );
  OAI22XL U3623 ( .A0(n782), .A1(n3907), .B0(n3104), .B1(n3920), .Y(n2022) );
  OAI22XL U3624 ( .A0(n783), .A1(n3907), .B0(n3103), .B1(n3921), .Y(n2023) );
  OAI22XL U3625 ( .A0(n784), .A1(n3907), .B0(n3102), .B1(n3921), .Y(n2024) );
  OAI22XL U3626 ( .A0(n785), .A1(n3907), .B0(n3089), .B1(n3921), .Y(n2025) );
  OAI22XL U3627 ( .A0(n786), .A1(n3907), .B0(n3101), .B1(n3921), .Y(n2026) );
  OAI22XL U3628 ( .A0(n787), .A1(n3908), .B0(n3100), .B1(n3921), .Y(n2027) );
  OAI22XL U3629 ( .A0(n788), .A1(n3908), .B0(n3099), .B1(n3921), .Y(n2028) );
  OAI22XL U3630 ( .A0(n789), .A1(n3908), .B0(n3098), .B1(n3921), .Y(n2029) );
  OAI22XL U3631 ( .A0(n790), .A1(n3908), .B0(n3088), .B1(n3921), .Y(n2030) );
  OAI22XL U3632 ( .A0(n791), .A1(n3908), .B0(n3152), .B1(n3921), .Y(n2031) );
  OAI22XL U3633 ( .A0(n792), .A1(n3908), .B0(n3151), .B1(n3921), .Y(n2032) );
  OAI22XL U3634 ( .A0(n793), .A1(n3908), .B0(n3168), .B1(n3921), .Y(n2033) );
  OAI22XL U3635 ( .A0(n794), .A1(n3908), .B0(n3170), .B1(n3922), .Y(n2034) );
  OAI22XL U3636 ( .A0(n795), .A1(n3908), .B0(n3159), .B1(n3922), .Y(n2035) );
  OAI22XL U3637 ( .A0(n796), .A1(n3908), .B0(n3150), .B1(n3922), .Y(n2036) );
  OAI22XL U3638 ( .A0(n797), .A1(n3908), .B0(n3161), .B1(n3922), .Y(n2037) );
  OAI22XL U3639 ( .A0(n798), .A1(n3908), .B0(n3149), .B1(n3922), .Y(n2038) );
  OAI22XL U3640 ( .A0(n799), .A1(n3909), .B0(n3163), .B1(n3922), .Y(n2039) );
  OAI22XL U3641 ( .A0(n800), .A1(n3909), .B0(n3165), .B1(n3922), .Y(n2040) );
  OAI22XL U3642 ( .A0(n801), .A1(n3909), .B0(n3167), .B1(n3922), .Y(n2041) );
  OAI22XL U3643 ( .A0(n802), .A1(n3909), .B0(n3169), .B1(n3922), .Y(n2042) );
  OAI22XL U3644 ( .A0(n803), .A1(n3909), .B0(n3148), .B1(n3922), .Y(n2043) );
  OAI22XL U3645 ( .A0(n804), .A1(n3909), .B0(n3147), .B1(n3922), .Y(n2044) );
  OAI22XL U3646 ( .A0(n805), .A1(n3909), .B0(n3158), .B1(n3923), .Y(n2045) );
  OAI22XL U3647 ( .A0(n806), .A1(n3909), .B0(n3157), .B1(n3923), .Y(n2046) );
  OAI22XL U3648 ( .A0(n807), .A1(n3909), .B0(n3166), .B1(n3923), .Y(n2047) );
  OAI22XL U3649 ( .A0(n808), .A1(n3909), .B0(n3156), .B1(n3923), .Y(n2048) );
  OAI22XL U3650 ( .A0(n809), .A1(n3909), .B0(n3160), .B1(n3923), .Y(n2049) );
  OAI22XL U3651 ( .A0(n810), .A1(n3909), .B0(n3162), .B1(n3923), .Y(n2050) );
  OAI22XL U3652 ( .A0(n811), .A1(n3910), .B0(n3164), .B1(n3923), .Y(n2051) );
  OAI22XL U3653 ( .A0(n812), .A1(n3910), .B0(n3155), .B1(n3923), .Y(n2052) );
  OAI22XL U3654 ( .A0(n813), .A1(n3910), .B0(n3154), .B1(n3923), .Y(n2053) );
  OAI22XL U3655 ( .A0(n814), .A1(n3910), .B0(n3153), .B1(n3923), .Y(n2054) );
  OAI22XL U3656 ( .A0(n815), .A1(n3910), .B0(n3097), .B1(n3923), .Y(n2055) );
  OAI22XL U3657 ( .A0(n816), .A1(n3910), .B0(n3093), .B1(n3924), .Y(n2056) );
  OAI22XL U3658 ( .A0(n817), .A1(n3910), .B0(n3092), .B1(n3924), .Y(n2057) );
  OAI22XL U3659 ( .A0(n818), .A1(n3910), .B0(n3091), .B1(n3924), .Y(n2058) );
  OAI22XL U3660 ( .A0(n819), .A1(n3910), .B0(n3090), .B1(n3924), .Y(n2059) );
  OAI22XL U3661 ( .A0(n820), .A1(n3910), .B0(n3096), .B1(n3924), .Y(n2060) );
  OAI22XL U3662 ( .A0(n821), .A1(n3910), .B0(n3095), .B1(n3924), .Y(n2061) );
  OAI22XL U3663 ( .A0(n822), .A1(n3910), .B0(n3094), .B1(n3924), .Y(n2062) );
  OAI22XL U3664 ( .A0(n823), .A1(n3911), .B0(n3179), .B1(n3924), .Y(n2063) );
  OAI22XL U3665 ( .A0(n824), .A1(n3911), .B0(n3178), .B1(n3924), .Y(n2064) );
  OAI22XL U3666 ( .A0(n825), .A1(n3911), .B0(n3177), .B1(n3924), .Y(n2065) );
  OAI22XL U3667 ( .A0(n826), .A1(n3911), .B0(n3176), .B1(n3924), .Y(n2066) );
  OAI22XL U3668 ( .A0(n827), .A1(n3911), .B0(n3187), .B1(n3925), .Y(n2067) );
  OAI22XL U3669 ( .A0(n828), .A1(n3911), .B0(n3186), .B1(n3925), .Y(n2068) );
  OAI22XL U3670 ( .A0(n829), .A1(n3911), .B0(n3185), .B1(n3925), .Y(n2069) );
  OAI22XL U3671 ( .A0(n830), .A1(n3911), .B0(n3184), .B1(n3925), .Y(n2070) );
  OAI22XL U3672 ( .A0(n831), .A1(n3911), .B0(n3183), .B1(n3925), .Y(n2071) );
  OAI22XL U3673 ( .A0(n832), .A1(n3911), .B0(n3182), .B1(n3925), .Y(n2072) );
  OAI22XL U3674 ( .A0(n833), .A1(n3911), .B0(n3146), .B1(n3925), .Y(n2073) );
  OAI22XL U3675 ( .A0(n834), .A1(n3911), .B0(n3145), .B1(n3925), .Y(n2074) );
  OAI22XL U3676 ( .A0(n835), .A1(n3912), .B0(n3144), .B1(n3925), .Y(n2075) );
  OAI22XL U3677 ( .A0(n836), .A1(n3912), .B0(n3143), .B1(n3925), .Y(n2076) );
  OAI22XL U3678 ( .A0(n837), .A1(n3912), .B0(n3142), .B1(n3925), .Y(n2077) );
  OAI22XL U3679 ( .A0(n838), .A1(n3912), .B0(n3139), .B1(n3926), .Y(n2078) );
  OAI22XL U3680 ( .A0(n839), .A1(n3912), .B0(n3138), .B1(n3926), .Y(n2079) );
  OAI22XL U3681 ( .A0(n840), .A1(n3912), .B0(n3137), .B1(n3926), .Y(n2080) );
  OAI22XL U3682 ( .A0(n841), .A1(n3912), .B0(n3136), .B1(n3926), .Y(n2081) );
  OAI22XL U3683 ( .A0(n842), .A1(n3912), .B0(n3141), .B1(n3926), .Y(n2082) );
  OAI22XL U3684 ( .A0(n843), .A1(n3912), .B0(n3135), .B1(n3926), .Y(n2083) );
  OAI22XL U3685 ( .A0(n844), .A1(n3912), .B0(n3140), .B1(n3926), .Y(n2084) );
  OAI22XL U3686 ( .A0(n845), .A1(n3912), .B0(n3172), .B1(n3926), .Y(n2085) );
  OAI22XL U3687 ( .A0(n846), .A1(n3912), .B0(n3180), .B1(n3926), .Y(n2086) );
  OAI22XL U3688 ( .A0(n847), .A1(n3913), .B0(n3173), .B1(n3926), .Y(n2087) );
  OAI22XL U3689 ( .A0(n848), .A1(n3913), .B0(n3171), .B1(n3926), .Y(n2088) );
  OAI22XL U3690 ( .A0(n849), .A1(n3913), .B0(n3189), .B1(n3917), .Y(n2089) );
  OAI22XL U3691 ( .A0(n850), .A1(n3913), .B0(n3188), .B1(n3928), .Y(n2090) );
  OAI22XL U3692 ( .A0(n851), .A1(n3913), .B0(n3175), .B1(n3918), .Y(n2091) );
  OAI22XL U3693 ( .A0(n852), .A1(n3913), .B0(n3181), .B1(n3919), .Y(n2092) );
  OAI22XL U3694 ( .A0(n853), .A1(n3913), .B0(n3174), .B1(n3922), .Y(n2093) );
  OAI22XL U3695 ( .A0(n882), .A1(n4101), .B0(n3080), .B1(n4114), .Y(n2122) );
  OAI22XL U3696 ( .A0(n884), .A1(n4101), .B0(n3081), .B1(n4114), .Y(n2124) );
  OAI22XL U3697 ( .A0(n885), .A1(n4101), .B0(n3079), .B1(n4114), .Y(n2125) );
  OAI22XL U3698 ( .A0(n886), .A1(n4101), .B0(n3078), .B1(n4114), .Y(n2126) );
  OAI22XL U3699 ( .A0(n887), .A1(n4101), .B0(n3077), .B1(n4115), .Y(n2127) );
  OAI22XL U3700 ( .A0(n888), .A1(n4101), .B0(n3076), .B1(n4115), .Y(n2128) );
  OAI22XL U3701 ( .A0(n889), .A1(n4102), .B0(n3086), .B1(n4115), .Y(n2129) );
  OAI22XL U3702 ( .A0(n890), .A1(n4102), .B0(n3085), .B1(n4115), .Y(n2130) );
  OAI22XL U3703 ( .A0(n891), .A1(n4102), .B0(n3084), .B1(n4115), .Y(n2131) );
  OAI22XL U3704 ( .A0(n892), .A1(n4102), .B0(n3083), .B1(n4115), .Y(n2132) );
  OAI22XL U3705 ( .A0(n893), .A1(n4102), .B0(n3082), .B1(n4115), .Y(n2133) );
  OAI22XL U3706 ( .A0(n894), .A1(n4102), .B0(n222), .B1(n4115), .Y(n2134) );
  OAI22XL U3707 ( .A0(n895), .A1(n4102), .B0(n223), .B1(n4115), .Y(n2135) );
  OAI22XL U3708 ( .A0(n896), .A1(n4102), .B0(n3130), .B1(n4115), .Y(n2136) );
  OAI22XL U3709 ( .A0(n897), .A1(n4102), .B0(n3129), .B1(n4115), .Y(n2137) );
  OAI22XL U3710 ( .A0(n898), .A1(n4102), .B0(n3128), .B1(n4116), .Y(n2138) );
  OAI22XL U3711 ( .A0(n899), .A1(n4102), .B0(n3127), .B1(n4116), .Y(n2139) );
  OAI22XL U3712 ( .A0(n900), .A1(n4102), .B0(n3126), .B1(n4116), .Y(n2140) );
  OAI22XL U3713 ( .A0(n901), .A1(n4103), .B0(n229), .B1(n4116), .Y(n2141) );
  OAI22XL U3714 ( .A0(n902), .A1(n4103), .B0(n3134), .B1(n4116), .Y(n2142) );
  OAI22XL U3715 ( .A0(n903), .A1(n4103), .B0(n3133), .B1(n4116), .Y(n2143) );
  OAI22XL U3716 ( .A0(n904), .A1(n4103), .B0(n3132), .B1(n4116), .Y(n2144) );
  OAI22XL U3717 ( .A0(n905), .A1(n4103), .B0(n3131), .B1(n4116), .Y(n2145) );
  OAI22XL U3718 ( .A0(n906), .A1(n4103), .B0(n3073), .B1(n4116), .Y(n2146) );
  OAI22XL U3719 ( .A0(n907), .A1(n4103), .B0(n3067), .B1(n4116), .Y(n2147) );
  OAI22XL U3720 ( .A0(n908), .A1(n4103), .B0(n3064), .B1(n4116), .Y(n2148) );
  OAI22XL U3721 ( .A0(n909), .A1(n4103), .B0(n3071), .B1(n4117), .Y(n2149) );
  OAI22XL U3722 ( .A0(n910), .A1(n4103), .B0(n3062), .B1(n4117), .Y(n2150) );
  OAI22XL U3723 ( .A0(n911), .A1(n4103), .B0(n3059), .B1(n4117), .Y(n2151) );
  OAI22XL U3724 ( .A0(n912), .A1(n4103), .B0(n3056), .B1(n4117), .Y(n2152) );
  OAI22XL U3725 ( .A0(n913), .A1(n4104), .B0(n3053), .B1(n4117), .Y(n2153) );
  OAI22XL U3726 ( .A0(n914), .A1(n4104), .B0(n242), .B1(n4117), .Y(n2154) );
  OAI22XL U3727 ( .A0(n915), .A1(n4104), .B0(n3125), .B1(n4117), .Y(n2155) );
  OAI22XL U3728 ( .A0(n916), .A1(n4104), .B0(n3124), .B1(n4117), .Y(n2156) );
  OAI22XL U3729 ( .A0(n917), .A1(n4104), .B0(n3123), .B1(n4117), .Y(n2157) );
  OAI22XL U3730 ( .A0(n918), .A1(n4104), .B0(n246), .B1(n4117), .Y(n2158) );
  OAI22XL U3731 ( .A0(n919), .A1(n4104), .B0(n3122), .B1(n4117), .Y(n2159) );
  OAI22XL U3732 ( .A0(n920), .A1(n4104), .B0(n3121), .B1(n4118), .Y(n2160) );
  OAI22XL U3733 ( .A0(n921), .A1(n4104), .B0(n3120), .B1(n4118), .Y(n2161) );
  OAI22XL U3734 ( .A0(n922), .A1(n4104), .B0(n3119), .B1(n4118), .Y(n2162) );
  OAI22XL U3735 ( .A0(n923), .A1(n4104), .B0(n3118), .B1(n4118), .Y(n2163) );
  OAI22XL U3736 ( .A0(n924), .A1(n4104), .B0(n3117), .B1(n4118), .Y(n2164) );
  OAI22XL U3737 ( .A0(n925), .A1(n4105), .B0(n3116), .B1(n4118), .Y(n2165) );
  OAI22XL U3738 ( .A0(n926), .A1(n4105), .B0(n3115), .B1(n4118), .Y(n2166) );
  OAI22XL U3739 ( .A0(n927), .A1(n4105), .B0(n3114), .B1(n4118), .Y(n2167) );
  OAI22XL U3740 ( .A0(n928), .A1(n4105), .B0(n3113), .B1(n4118), .Y(n2168) );
  OAI22XL U3741 ( .A0(n929), .A1(n4105), .B0(n3112), .B1(n4118), .Y(n2169) );
  OAI22XL U3742 ( .A0(n930), .A1(n4105), .B0(n3111), .B1(n4118), .Y(n2170) );
  OAI22XL U3743 ( .A0(n931), .A1(n4105), .B0(n3110), .B1(n4119), .Y(n2171) );
  OAI22XL U3744 ( .A0(n932), .A1(n4105), .B0(n3109), .B1(n4119), .Y(n2172) );
  OAI22XL U3745 ( .A0(n933), .A1(n4105), .B0(n3108), .B1(n4119), .Y(n2173) );
  OAI22XL U3746 ( .A0(n934), .A1(n4105), .B0(n3107), .B1(n4119), .Y(n2174) );
  OAI22XL U3747 ( .A0(n935), .A1(n4105), .B0(n3106), .B1(n4119), .Y(n2175) );
  OAI22XL U3748 ( .A0(n936), .A1(n4105), .B0(n3105), .B1(n4119), .Y(n2176) );
  OAI22XL U3749 ( .A0(n937), .A1(n4106), .B0(n3104), .B1(n4119), .Y(n2177) );
  OAI22XL U3750 ( .A0(n938), .A1(n4106), .B0(n3103), .B1(n4119), .Y(n2178) );
  OAI22XL U3751 ( .A0(n939), .A1(n4106), .B0(n3102), .B1(n4119), .Y(n2179) );
  OAI22XL U3752 ( .A0(n940), .A1(n4106), .B0(n3089), .B1(n4119), .Y(n2180) );
  OAI22XL U3753 ( .A0(n941), .A1(n4106), .B0(n3101), .B1(n4119), .Y(n2181) );
  OAI22XL U3754 ( .A0(n942), .A1(n4106), .B0(n3100), .B1(n4120), .Y(n2182) );
  OAI22XL U3755 ( .A0(n943), .A1(n4106), .B0(n3099), .B1(n4120), .Y(n2183) );
  OAI22XL U3756 ( .A0(n944), .A1(n4106), .B0(n3098), .B1(n4120), .Y(n2184) );
  OAI22XL U3757 ( .A0(n945), .A1(n4106), .B0(n3088), .B1(n4120), .Y(n2185) );
  OAI22XL U3758 ( .A0(n946), .A1(n4106), .B0(n3152), .B1(n4120), .Y(n2186) );
  OAI22XL U3759 ( .A0(n947), .A1(n4106), .B0(n3151), .B1(n4120), .Y(n2187) );
  OAI22XL U3760 ( .A0(n948), .A1(n4106), .B0(n3168), .B1(n4120), .Y(n2188) );
  OAI22XL U3761 ( .A0(n949), .A1(n4107), .B0(n3170), .B1(n4120), .Y(n2189) );
  OAI22XL U3762 ( .A0(n950), .A1(n4107), .B0(n3159), .B1(n4120), .Y(n2190) );
  OAI22XL U3763 ( .A0(n951), .A1(n4107), .B0(n3150), .B1(n4120), .Y(n2191) );
  OAI22XL U3764 ( .A0(n952), .A1(n4107), .B0(n3161), .B1(n4120), .Y(n2192) );
  OAI22XL U3765 ( .A0(n953), .A1(n4107), .B0(n3149), .B1(n4121), .Y(n2193) );
  OAI22XL U3766 ( .A0(n954), .A1(n4107), .B0(n3163), .B1(n4121), .Y(n2194) );
  OAI22XL U3767 ( .A0(n955), .A1(n4107), .B0(n3165), .B1(n4121), .Y(n2195) );
  OAI22XL U3768 ( .A0(n956), .A1(n4107), .B0(n3167), .B1(n4121), .Y(n2196) );
  OAI22XL U3769 ( .A0(n957), .A1(n4107), .B0(n3169), .B1(n4121), .Y(n2197) );
  OAI22XL U3770 ( .A0(n958), .A1(n4107), .B0(n3148), .B1(n4121), .Y(n2198) );
  OAI22XL U3771 ( .A0(n959), .A1(n4107), .B0(n3147), .B1(n4121), .Y(n2199) );
  OAI22XL U3772 ( .A0(n960), .A1(n4107), .B0(n3158), .B1(n4121), .Y(n2200) );
  OAI22XL U3773 ( .A0(n961), .A1(n4108), .B0(n3157), .B1(n4121), .Y(n2201) );
  OAI22XL U3774 ( .A0(n962), .A1(n4108), .B0(n3166), .B1(n4121), .Y(n2202) );
  OAI22XL U3775 ( .A0(n963), .A1(n4108), .B0(n3156), .B1(n4121), .Y(n2203) );
  OAI22XL U3776 ( .A0(n964), .A1(n4108), .B0(n3160), .B1(n4122), .Y(n2204) );
  OAI22XL U3777 ( .A0(n965), .A1(n4108), .B0(n3162), .B1(n4122), .Y(n2205) );
  OAI22XL U3778 ( .A0(n966), .A1(n4108), .B0(n3164), .B1(n4122), .Y(n2206) );
  OAI22XL U3779 ( .A0(n967), .A1(n4108), .B0(n3155), .B1(n4122), .Y(n2207) );
  OAI22XL U3780 ( .A0(n968), .A1(n4108), .B0(n3154), .B1(n4122), .Y(n2208) );
  OAI22XL U3781 ( .A0(n969), .A1(n4108), .B0(n3153), .B1(n4122), .Y(n2209) );
  OAI22XL U3782 ( .A0(n970), .A1(n4108), .B0(n3097), .B1(n4122), .Y(n2210) );
  OAI22XL U3783 ( .A0(n971), .A1(n4108), .B0(n3093), .B1(n4122), .Y(n2211) );
  OAI22XL U3784 ( .A0(n972), .A1(n4108), .B0(n3092), .B1(n4122), .Y(n2212) );
  OAI22XL U3785 ( .A0(n973), .A1(n4109), .B0(n3091), .B1(n4122), .Y(n2213) );
  OAI22XL U3786 ( .A0(n974), .A1(n4109), .B0(n3090), .B1(n4122), .Y(n2214) );
  OAI22XL U3787 ( .A0(n975), .A1(n4109), .B0(n3096), .B1(n4123), .Y(n2215) );
  OAI22XL U3788 ( .A0(n976), .A1(n4109), .B0(n3095), .B1(n4123), .Y(n2216) );
  OAI22XL U3789 ( .A0(n977), .A1(n4109), .B0(n3094), .B1(n4123), .Y(n2217) );
  OAI22XL U3790 ( .A0(n978), .A1(n4109), .B0(n3179), .B1(n4123), .Y(n2218) );
  OAI22XL U3791 ( .A0(n979), .A1(n4109), .B0(n3178), .B1(n4123), .Y(n2219) );
  OAI22XL U3792 ( .A0(n980), .A1(n4109), .B0(n3177), .B1(n4123), .Y(n2220) );
  OAI22XL U3793 ( .A0(n981), .A1(n4109), .B0(n3176), .B1(n4123), .Y(n2221) );
  OAI22XL U3794 ( .A0(n982), .A1(n4109), .B0(n3187), .B1(n4123), .Y(n2222) );
  OAI22XL U3795 ( .A0(n983), .A1(n4109), .B0(n3186), .B1(n4123), .Y(n2223) );
  OAI22XL U3796 ( .A0(n984), .A1(n4109), .B0(n3185), .B1(n4123), .Y(n2224) );
  OAI22XL U3797 ( .A0(n985), .A1(n4110), .B0(n3184), .B1(n4123), .Y(n2225) );
  OAI22XL U3798 ( .A0(n986), .A1(n4110), .B0(n3183), .B1(n4124), .Y(n2226) );
  OAI22XL U3799 ( .A0(n987), .A1(n4110), .B0(n3182), .B1(n4124), .Y(n2227) );
  OAI22XL U3800 ( .A0(n988), .A1(n4110), .B0(n3146), .B1(n4124), .Y(n2228) );
  OAI22XL U3801 ( .A0(n989), .A1(n4110), .B0(n3145), .B1(n4124), .Y(n2229) );
  OAI22XL U3802 ( .A0(n990), .A1(n4110), .B0(n3144), .B1(n4124), .Y(n2230) );
  OAI22XL U3803 ( .A0(n991), .A1(n4110), .B0(n3143), .B1(n4124), .Y(n2231) );
  OAI22XL U3804 ( .A0(n992), .A1(n4110), .B0(n3142), .B1(n4124), .Y(n2232) );
  OAI22XL U3805 ( .A0(n993), .A1(n4110), .B0(n3139), .B1(n4124), .Y(n2233) );
  OAI22XL U3806 ( .A0(n994), .A1(n4110), .B0(n3138), .B1(n4124), .Y(n2234) );
  OAI22XL U3807 ( .A0(n995), .A1(n4110), .B0(n3137), .B1(n4124), .Y(n2235) );
  OAI22XL U3808 ( .A0(n996), .A1(n4110), .B0(n3136), .B1(n4124), .Y(n2236) );
  OAI22XL U3809 ( .A0(n997), .A1(n4104), .B0(n3141), .B1(n4123), .Y(n2237) );
  OAI22XL U3810 ( .A0(n998), .A1(n4104), .B0(n3135), .B1(n4124), .Y(n2238) );
  OAI22XL U3811 ( .A0(n999), .A1(n4104), .B0(n3140), .B1(n4123), .Y(n2239) );
  OAI22XL U3812 ( .A0(n1000), .A1(n4104), .B0(n3172), .B1(n4124), .Y(n2240) );
  OAI22XL U3813 ( .A0(n1001), .A1(n4104), .B0(n3180), .B1(n4123), .Y(n2241) );
  OAI22XL U3814 ( .A0(n1002), .A1(n4102), .B0(n3173), .B1(n4124), .Y(n2242) );
  OAI22XL U3815 ( .A0(n1003), .A1(n4101), .B0(n3171), .B1(n4118), .Y(n2243) );
  OAI22XL U3816 ( .A0(n1004), .A1(n4102), .B0(n3189), .B1(n4117), .Y(n2244) );
  OAI22XL U3817 ( .A0(n1005), .A1(n4104), .B0(n3188), .B1(n4115), .Y(n2245) );
  OAI22XL U3818 ( .A0(n1006), .A1(n4101), .B0(n3175), .B1(n4119), .Y(n2246) );
  OAI22XL U3819 ( .A0(n1007), .A1(n4104), .B0(n3181), .B1(n4123), .Y(n2247) );
  OAI22XL U3820 ( .A0(n1008), .A1(n4099), .B0(n3174), .B1(n4111), .Y(n2248) );
  OAI22XL U3821 ( .A0(n1037), .A1(n4071), .B0(n3080), .B1(n4096), .Y(n2277) );
  OAI22XL U3822 ( .A0(n1038), .A1(n4071), .B0(n211), .B1(n4094), .Y(n2278) );
  OAI22XL U3823 ( .A0(n1039), .A1(n4071), .B0(n3081), .B1(n4085), .Y(n2279) );
  OAI22XL U3824 ( .A0(n1040), .A1(n4071), .B0(n3079), .B1(n4095), .Y(n2280) );
  OAI22XL U3825 ( .A0(n1041), .A1(n4071), .B0(n3078), .B1(n4084), .Y(n2281) );
  OAI22XL U3826 ( .A0(n1042), .A1(n4071), .B0(n3077), .B1(n4084), .Y(n2282) );
  OAI22XL U3827 ( .A0(n1043), .A1(n4071), .B0(n3076), .B1(n4084), .Y(n2283) );
  OAI22XL U3828 ( .A0(n1044), .A1(n4071), .B0(n3086), .B1(n4084), .Y(n2284) );
  OAI22XL U3829 ( .A0(n1045), .A1(n4071), .B0(n3085), .B1(n4084), .Y(n2285) );
  OAI22XL U3830 ( .A0(n1046), .A1(n4071), .B0(n3084), .B1(n4084), .Y(n2286) );
  OAI22XL U3831 ( .A0(n1047), .A1(n4071), .B0(n3083), .B1(n4084), .Y(n2287) );
  OAI22XL U3832 ( .A0(n1048), .A1(n4071), .B0(n3082), .B1(n4084), .Y(n2288) );
  OAI22XL U3833 ( .A0(n1049), .A1(n4072), .B0(n222), .B1(n4085), .Y(n2289) );
  OAI22XL U3834 ( .A0(n1050), .A1(n4072), .B0(n223), .B1(n4085), .Y(n2290) );
  OAI22XL U3835 ( .A0(n1051), .A1(n4072), .B0(n3130), .B1(n4085), .Y(n2291) );
  OAI22XL U3836 ( .A0(n1052), .A1(n4072), .B0(n3129), .B1(n4085), .Y(n2292) );
  OAI22XL U3837 ( .A0(n1053), .A1(n4072), .B0(n3128), .B1(n4085), .Y(n2293) );
  OAI22XL U3838 ( .A0(n1054), .A1(n4072), .B0(n3127), .B1(n4085), .Y(n2294) );
  OAI22XL U3839 ( .A0(n1055), .A1(n4072), .B0(n3126), .B1(n4085), .Y(n2295) );
  OAI22XL U3840 ( .A0(n1056), .A1(n4072), .B0(n229), .B1(n4085), .Y(n2296) );
  OAI22XL U3841 ( .A0(n1057), .A1(n4072), .B0(n3134), .B1(n4085), .Y(n2297) );
  OAI22XL U3842 ( .A0(n1058), .A1(n4072), .B0(n3133), .B1(n4085), .Y(n2298) );
  OAI22XL U3843 ( .A0(n1059), .A1(n4072), .B0(n3132), .B1(n4085), .Y(n2299) );
  OAI22XL U3844 ( .A0(n1060), .A1(n4072), .B0(n3131), .B1(n4086), .Y(n2300) );
  OAI22XL U3845 ( .A0(n1061), .A1(n4073), .B0(n3074), .B1(n4086), .Y(n2301) );
  OAI22XL U3846 ( .A0(n1062), .A1(n4073), .B0(n3068), .B1(n4086), .Y(n2302) );
  OAI22XL U3847 ( .A0(n1063), .A1(n4073), .B0(n3065), .B1(n4086), .Y(n2303) );
  OAI22XL U3848 ( .A0(n1064), .A1(n4073), .B0(n3071), .B1(n4086), .Y(n2304) );
  OAI22XL U3849 ( .A0(n1065), .A1(n4073), .B0(n3062), .B1(n4086), .Y(n2305) );
  OAI22XL U3850 ( .A0(n1066), .A1(n4073), .B0(n3059), .B1(n4086), .Y(n2306) );
  OAI22XL U3851 ( .A0(n1067), .A1(n4073), .B0(n3056), .B1(n4086), .Y(n2307) );
  OAI22XL U3852 ( .A0(n1068), .A1(n4073), .B0(n3053), .B1(n4086), .Y(n2308) );
  OAI22XL U3853 ( .A0(n1069), .A1(n4073), .B0(n242), .B1(n4086), .Y(n2309) );
  OAI22XL U3854 ( .A0(n1070), .A1(n4073), .B0(n3125), .B1(n4086), .Y(n2310) );
  OAI22XL U3855 ( .A0(n1071), .A1(n4073), .B0(n3124), .B1(n4087), .Y(n2311) );
  OAI22XL U3856 ( .A0(n1072), .A1(n4073), .B0(n3123), .B1(n4087), .Y(n2312) );
  OAI22XL U3857 ( .A0(n1073), .A1(n4074), .B0(n246), .B1(n4087), .Y(n2313) );
  OAI22XL U3858 ( .A0(n1074), .A1(n4074), .B0(n3122), .B1(n4087), .Y(n2314) );
  OAI22XL U3859 ( .A0(n1075), .A1(n4074), .B0(n3121), .B1(n4087), .Y(n2315) );
  OAI22XL U3860 ( .A0(n1076), .A1(n4074), .B0(n3120), .B1(n4087), .Y(n2316) );
  OAI22XL U3861 ( .A0(n1077), .A1(n4074), .B0(n3119), .B1(n4087), .Y(n2317) );
  OAI22XL U3862 ( .A0(n1078), .A1(n4074), .B0(n3118), .B1(n4087), .Y(n2318) );
  OAI22XL U3863 ( .A0(n1079), .A1(n4074), .B0(n3117), .B1(n4087), .Y(n2319) );
  OAI22XL U3864 ( .A0(n1080), .A1(n4074), .B0(n3116), .B1(n4087), .Y(n2320) );
  OAI22XL U3865 ( .A0(n1081), .A1(n4074), .B0(n3115), .B1(n4087), .Y(n2321) );
  OAI22XL U3866 ( .A0(n1082), .A1(n4074), .B0(n3114), .B1(n4088), .Y(n2322) );
  OAI22XL U3867 ( .A0(n1083), .A1(n4074), .B0(n3113), .B1(n4088), .Y(n2323) );
  OAI22XL U3868 ( .A0(n1084), .A1(n4074), .B0(n3112), .B1(n4088), .Y(n2324) );
  OAI22XL U3869 ( .A0(n1085), .A1(n4075), .B0(n3111), .B1(n4088), .Y(n2325) );
  OAI22XL U3870 ( .A0(n1086), .A1(n4075), .B0(n3110), .B1(n4088), .Y(n2326) );
  OAI22XL U3871 ( .A0(n1087), .A1(n4075), .B0(n3109), .B1(n4088), .Y(n2327) );
  OAI22XL U3872 ( .A0(n1088), .A1(n4075), .B0(n3108), .B1(n4088), .Y(n2328) );
  OAI22XL U3873 ( .A0(n1089), .A1(n4075), .B0(n3107), .B1(n4088), .Y(n2329) );
  OAI22XL U3874 ( .A0(n1090), .A1(n4075), .B0(n3106), .B1(n4088), .Y(n2330) );
  OAI22XL U3875 ( .A0(n1091), .A1(n4075), .B0(n3105), .B1(n4088), .Y(n2331) );
  OAI22XL U3876 ( .A0(n1092), .A1(n4075), .B0(n3104), .B1(n4088), .Y(n2332) );
  OAI22XL U3877 ( .A0(n1093), .A1(n4075), .B0(n3103), .B1(n4089), .Y(n2333) );
  OAI22XL U3878 ( .A0(n1094), .A1(n4075), .B0(n3102), .B1(n4089), .Y(n2334) );
  OAI22XL U3879 ( .A0(n1095), .A1(n4075), .B0(n3089), .B1(n4089), .Y(n2335) );
  OAI22XL U3880 ( .A0(n1096), .A1(n4075), .B0(n3101), .B1(n4089), .Y(n2336) );
  OAI22XL U3881 ( .A0(n1097), .A1(n4076), .B0(n3100), .B1(n4089), .Y(n2337) );
  OAI22XL U3882 ( .A0(n1098), .A1(n4076), .B0(n3099), .B1(n4089), .Y(n2338) );
  OAI22XL U3883 ( .A0(n1099), .A1(n4076), .B0(n3098), .B1(n4089), .Y(n2339) );
  OAI22XL U3884 ( .A0(n1100), .A1(n4076), .B0(n3088), .B1(n4089), .Y(n2340) );
  OAI22XL U3885 ( .A0(n1101), .A1(n4076), .B0(n3152), .B1(n4089), .Y(n2341) );
  OAI22XL U3886 ( .A0(n1102), .A1(n4076), .B0(n3151), .B1(n4089), .Y(n2342) );
  OAI22XL U3887 ( .A0(n1103), .A1(n4076), .B0(n3168), .B1(n4089), .Y(n2343) );
  OAI22XL U3888 ( .A0(n1104), .A1(n4076), .B0(n3170), .B1(n4090), .Y(n2344) );
  OAI22XL U3889 ( .A0(n1105), .A1(n4076), .B0(n3159), .B1(n4090), .Y(n2345) );
  OAI22XL U3890 ( .A0(n1106), .A1(n4076), .B0(n3150), .B1(n4090), .Y(n2346) );
  OAI22XL U3891 ( .A0(n1107), .A1(n4076), .B0(n3161), .B1(n4090), .Y(n2347) );
  OAI22XL U3892 ( .A0(n1108), .A1(n4076), .B0(n3149), .B1(n4090), .Y(n2348) );
  OAI22XL U3893 ( .A0(n1109), .A1(n4077), .B0(n3163), .B1(n4090), .Y(n2349) );
  OAI22XL U3894 ( .A0(n1110), .A1(n4077), .B0(n3165), .B1(n4090), .Y(n2350) );
  OAI22XL U3895 ( .A0(n1111), .A1(n4077), .B0(n3167), .B1(n4090), .Y(n2351) );
  OAI22XL U3896 ( .A0(n1112), .A1(n4077), .B0(n3169), .B1(n4090), .Y(n2352) );
  OAI22XL U3897 ( .A0(n1113), .A1(n4077), .B0(n3148), .B1(n4090), .Y(n2353) );
  OAI22XL U3898 ( .A0(n1114), .A1(n4077), .B0(n3147), .B1(n4090), .Y(n2354) );
  OAI22XL U3899 ( .A0(n1115), .A1(n4077), .B0(n3158), .B1(n4091), .Y(n2355) );
  OAI22XL U3900 ( .A0(n1116), .A1(n4077), .B0(n3157), .B1(n4091), .Y(n2356) );
  OAI22XL U3901 ( .A0(n1117), .A1(n4077), .B0(n3166), .B1(n4091), .Y(n2357) );
  OAI22XL U3902 ( .A0(n1118), .A1(n4077), .B0(n3156), .B1(n4091), .Y(n2358) );
  OAI22XL U3903 ( .A0(n1119), .A1(n4077), .B0(n3160), .B1(n4091), .Y(n2359) );
  OAI22XL U3904 ( .A0(n1120), .A1(n4077), .B0(n3162), .B1(n4091), .Y(n2360) );
  OAI22XL U3905 ( .A0(n1121), .A1(n4078), .B0(n3164), .B1(n4091), .Y(n2361) );
  OAI22XL U3906 ( .A0(n1122), .A1(n4078), .B0(n3155), .B1(n4091), .Y(n2362) );
  OAI22XL U3907 ( .A0(n1123), .A1(n4078), .B0(n3154), .B1(n4091), .Y(n2363) );
  OAI22XL U3908 ( .A0(n1124), .A1(n4078), .B0(n3153), .B1(n4091), .Y(n2364) );
  OAI22XL U3909 ( .A0(n1125), .A1(n4078), .B0(n3097), .B1(n4091), .Y(n2365) );
  OAI22XL U3910 ( .A0(n1126), .A1(n4078), .B0(n3093), .B1(n4092), .Y(n2366) );
  OAI22XL U3911 ( .A0(n1127), .A1(n4078), .B0(n3092), .B1(n4092), .Y(n2367) );
  OAI22XL U3912 ( .A0(n1128), .A1(n4078), .B0(n3091), .B1(n4092), .Y(n2368) );
  OAI22XL U3913 ( .A0(n1129), .A1(n4078), .B0(n3090), .B1(n4092), .Y(n2369) );
  OAI22XL U3914 ( .A0(n1130), .A1(n4078), .B0(n3096), .B1(n4092), .Y(n2370) );
  OAI22XL U3915 ( .A0(n1131), .A1(n4078), .B0(n3095), .B1(n4092), .Y(n2371) );
  OAI22XL U3916 ( .A0(n1132), .A1(n4078), .B0(n3094), .B1(n4092), .Y(n2372) );
  OAI22XL U3917 ( .A0(n1133), .A1(n4079), .B0(n3179), .B1(n4092), .Y(n2373) );
  OAI22XL U3918 ( .A0(n1134), .A1(n4079), .B0(n3178), .B1(n4092), .Y(n2374) );
  OAI22XL U3919 ( .A0(n1135), .A1(n4079), .B0(n3177), .B1(n4092), .Y(n2375) );
  OAI22XL U3920 ( .A0(n1136), .A1(n4079), .B0(n3176), .B1(n4092), .Y(n2376) );
  OAI22XL U3921 ( .A0(n1137), .A1(n4079), .B0(n3187), .B1(n4093), .Y(n2377) );
  OAI22XL U3922 ( .A0(n1138), .A1(n4079), .B0(n3186), .B1(n4093), .Y(n2378) );
  OAI22XL U3923 ( .A0(n1139), .A1(n4079), .B0(n3185), .B1(n4093), .Y(n2379) );
  OAI22XL U3924 ( .A0(n1140), .A1(n4079), .B0(n3184), .B1(n4093), .Y(n2380) );
  OAI22XL U3925 ( .A0(n1141), .A1(n4079), .B0(n3183), .B1(n4093), .Y(n2381) );
  OAI22XL U3926 ( .A0(n1142), .A1(n4079), .B0(n3182), .B1(n4093), .Y(n2382) );
  OAI22XL U3927 ( .A0(n1143), .A1(n4079), .B0(n3146), .B1(n4093), .Y(n2383) );
  OAI22XL U3928 ( .A0(n1144), .A1(n4079), .B0(n3145), .B1(n4093), .Y(n2384) );
  OAI22XL U3929 ( .A0(n1145), .A1(n4080), .B0(n3144), .B1(n4093), .Y(n2385) );
  OAI22XL U3930 ( .A0(n1146), .A1(n4080), .B0(n3143), .B1(n4093), .Y(n2386) );
  OAI22XL U3931 ( .A0(n1147), .A1(n4080), .B0(n3142), .B1(n4093), .Y(n2387) );
  OAI22XL U3932 ( .A0(n1148), .A1(n4080), .B0(n3139), .B1(n4094), .Y(n2388) );
  OAI22XL U3933 ( .A0(n1149), .A1(n4080), .B0(n3138), .B1(n4094), .Y(n2389) );
  OAI22XL U3934 ( .A0(n1150), .A1(n4080), .B0(n3137), .B1(n4094), .Y(n2390) );
  OAI22XL U3935 ( .A0(n1151), .A1(n4080), .B0(n3136), .B1(n4094), .Y(n2391) );
  OAI22XL U3936 ( .A0(n1152), .A1(n4080), .B0(n3141), .B1(n4094), .Y(n2392) );
  OAI22XL U3937 ( .A0(n1153), .A1(n4080), .B0(n3135), .B1(n4094), .Y(n2393) );
  OAI22XL U3938 ( .A0(n1154), .A1(n4080), .B0(n3140), .B1(n4094), .Y(n2394) );
  OAI22XL U3939 ( .A0(n1155), .A1(n4080), .B0(n3172), .B1(n4094), .Y(n2395) );
  OAI22XL U3940 ( .A0(n1156), .A1(n4080), .B0(n3180), .B1(n4094), .Y(n2396) );
  OAI22XL U3941 ( .A0(n1157), .A1(n4081), .B0(n3173), .B1(n4094), .Y(n2397) );
  OAI22XL U3942 ( .A0(n1158), .A1(n4081), .B0(n3171), .B1(n4094), .Y(n2398) );
  OAI22XL U3943 ( .A0(n1159), .A1(n4081), .B0(n3189), .B1(n4085), .Y(n2399) );
  OAI22XL U3944 ( .A0(n1160), .A1(n4081), .B0(n3188), .B1(n4096), .Y(n2400) );
  OAI22XL U3945 ( .A0(n1161), .A1(n4081), .B0(n3175), .B1(n4086), .Y(n2401) );
  OAI22XL U3946 ( .A0(n1162), .A1(n4081), .B0(n3181), .B1(n4087), .Y(n2402) );
  OAI22XL U3947 ( .A0(n1163), .A1(n4081), .B0(n3174), .B1(n4090), .Y(n2403) );
  OAI22XL U3948 ( .A0(n1192), .A1(n4043), .B0(n3080), .B1(n4068), .Y(n2432) );
  OAI22XL U3949 ( .A0(n1193), .A1(n4043), .B0(n211), .B1(n4055), .Y(n2433) );
  OAI22XL U3950 ( .A0(n1194), .A1(n4043), .B0(n3081), .B1(n4065), .Y(n2434) );
  OAI22XL U3951 ( .A0(n1195), .A1(n4043), .B0(n3079), .B1(n4067), .Y(n2435) );
  OAI22XL U3952 ( .A0(n1196), .A1(n4043), .B0(n3078), .B1(n4060), .Y(n2436) );
  OAI22XL U3953 ( .A0(n1197), .A1(n4043), .B0(n3077), .B1(n4063), .Y(n2437) );
  OAI22XL U3954 ( .A0(n1198), .A1(n4043), .B0(n3076), .B1(n4059), .Y(n2438) );
  OAI22XL U3955 ( .A0(n1199), .A1(n4043), .B0(n3086), .B1(n4060), .Y(n2439) );
  OAI22XL U3956 ( .A0(n1200), .A1(n4043), .B0(n3085), .B1(n4063), .Y(n2440) );
  OAI22XL U3957 ( .A0(n1201), .A1(n4043), .B0(n3084), .B1(n4059), .Y(n2441) );
  OAI22XL U3958 ( .A0(n1202), .A1(n4043), .B0(n3083), .B1(n4067), .Y(n2442) );
  OAI22XL U3959 ( .A0(n1203), .A1(n4043), .B0(n3082), .B1(n4068), .Y(n2443) );
  OAI22XL U3960 ( .A0(n1204), .A1(n4044), .B0(n222), .B1(n4056), .Y(n2444) );
  OAI22XL U3961 ( .A0(n1205), .A1(n4044), .B0(n223), .B1(n4056), .Y(n2445) );
  OAI22XL U3962 ( .A0(n1206), .A1(n4044), .B0(n3130), .B1(n4056), .Y(n2446) );
  OAI22XL U3963 ( .A0(n1207), .A1(n4044), .B0(n3129), .B1(n4056), .Y(n2447) );
  OAI22XL U3964 ( .A0(n1208), .A1(n4044), .B0(n3128), .B1(n4056), .Y(n2448) );
  OAI22XL U3965 ( .A0(n1209), .A1(n4044), .B0(n3127), .B1(n4056), .Y(n2449) );
  OAI22XL U3966 ( .A0(n1210), .A1(n4044), .B0(n3126), .B1(n4056), .Y(n2450) );
  OAI22XL U3967 ( .A0(n1211), .A1(n4044), .B0(n229), .B1(n4056), .Y(n2451) );
  OAI22XL U3968 ( .A0(n1212), .A1(n4044), .B0(n3134), .B1(n4056), .Y(n2452) );
  OAI22XL U3969 ( .A0(n1213), .A1(n4044), .B0(n3133), .B1(n4056), .Y(n2453) );
  OAI22XL U3970 ( .A0(n1214), .A1(n4044), .B0(n3132), .B1(n4056), .Y(n2454) );
  OAI22XL U3971 ( .A0(n1215), .A1(n4044), .B0(n3131), .B1(n4057), .Y(n2455) );
  OAI22XL U3972 ( .A0(n1216), .A1(n4045), .B0(n3073), .B1(n4057), .Y(n2456) );
  OAI22XL U3973 ( .A0(n1217), .A1(n4045), .B0(n3067), .B1(n4057), .Y(n2457) );
  OAI22XL U3974 ( .A0(n1218), .A1(n4045), .B0(n3064), .B1(n4057), .Y(n2458) );
  OAI22XL U3975 ( .A0(n1219), .A1(n4045), .B0(n3070), .B1(n4057), .Y(n2459) );
  OAI22XL U3976 ( .A0(n1220), .A1(n4045), .B0(n3061), .B1(n4057), .Y(n2460) );
  OAI22XL U3977 ( .A0(n1221), .A1(n4045), .B0(n3058), .B1(n4057), .Y(n2461) );
  OAI22XL U3978 ( .A0(n1222), .A1(n4045), .B0(n3055), .B1(n4057), .Y(n2462) );
  OAI22XL U3979 ( .A0(n1223), .A1(n4045), .B0(n3053), .B1(n4057), .Y(n2463) );
  OAI22XL U3980 ( .A0(n1224), .A1(n4045), .B0(n242), .B1(n4057), .Y(n2464) );
  OAI22XL U3981 ( .A0(n1225), .A1(n4045), .B0(n3125), .B1(n4057), .Y(n2465) );
  OAI22XL U3982 ( .A0(n1226), .A1(n4045), .B0(n3124), .B1(n4058), .Y(n2466) );
  OAI22XL U3983 ( .A0(n1227), .A1(n4045), .B0(n3123), .B1(n4058), .Y(n2467) );
  OAI22XL U3984 ( .A0(n1228), .A1(n4046), .B0(n246), .B1(n4058), .Y(n2468) );
  OAI22XL U3985 ( .A0(n1229), .A1(n4046), .B0(n3122), .B1(n4058), .Y(n2469) );
  OAI22XL U3986 ( .A0(n1230), .A1(n4046), .B0(n3121), .B1(n4058), .Y(n2470) );
  OAI22XL U3987 ( .A0(n1231), .A1(n4046), .B0(n3120), .B1(n4058), .Y(n2471) );
  OAI22XL U3988 ( .A0(n1232), .A1(n4046), .B0(n3119), .B1(n4058), .Y(n2472) );
  OAI22XL U3989 ( .A0(n1233), .A1(n4046), .B0(n3118), .B1(n4058), .Y(n2473) );
  OAI22XL U3990 ( .A0(n1234), .A1(n4046), .B0(n3117), .B1(n4058), .Y(n2474) );
  OAI22XL U3991 ( .A0(n1235), .A1(n4046), .B0(n3116), .B1(n4058), .Y(n2475) );
  OAI22XL U3992 ( .A0(n1236), .A1(n4046), .B0(n3115), .B1(n4058), .Y(n2476) );
  OAI22XL U3993 ( .A0(n1237), .A1(n4046), .B0(n3114), .B1(n4059), .Y(n2477) );
  OAI22XL U3994 ( .A0(n1238), .A1(n4046), .B0(n3113), .B1(n4059), .Y(n2478) );
  OAI22XL U3995 ( .A0(n1239), .A1(n4046), .B0(n3112), .B1(n4059), .Y(n2479) );
  OAI22XL U3996 ( .A0(n1240), .A1(n4047), .B0(n3111), .B1(n4059), .Y(n2480) );
  OAI22XL U3997 ( .A0(n1241), .A1(n4047), .B0(n3110), .B1(n4059), .Y(n2481) );
  OAI22XL U3998 ( .A0(n1242), .A1(n4047), .B0(n3109), .B1(n4059), .Y(n2482) );
  OAI22XL U3999 ( .A0(n1243), .A1(n4047), .B0(n3108), .B1(n4059), .Y(n2483) );
  OAI22XL U4000 ( .A0(n1244), .A1(n4047), .B0(n3107), .B1(n4059), .Y(n2484) );
  OAI22XL U4001 ( .A0(n1245), .A1(n4047), .B0(n3106), .B1(n4059), .Y(n2485) );
  OAI22XL U4002 ( .A0(n1246), .A1(n4047), .B0(n3105), .B1(n4059), .Y(n2486) );
  OAI22XL U4003 ( .A0(n1247), .A1(n4047), .B0(n3104), .B1(n4059), .Y(n2487) );
  OAI22XL U4004 ( .A0(n1248), .A1(n4047), .B0(n3103), .B1(n4060), .Y(n2488) );
  OAI22XL U4005 ( .A0(n1249), .A1(n4047), .B0(n3102), .B1(n4060), .Y(n2489) );
  OAI22XL U4006 ( .A0(n1250), .A1(n4047), .B0(n3089), .B1(n4060), .Y(n2490) );
  OAI22XL U4007 ( .A0(n1251), .A1(n4047), .B0(n3101), .B1(n4060), .Y(n2491) );
  OAI22XL U4008 ( .A0(n1252), .A1(n4048), .B0(n3100), .B1(n4060), .Y(n2492) );
  OAI22XL U4009 ( .A0(n1253), .A1(n4048), .B0(n3099), .B1(n4060), .Y(n2493) );
  OAI22XL U4010 ( .A0(n1254), .A1(n4048), .B0(n3098), .B1(n4060), .Y(n2494) );
  OAI22XL U4011 ( .A0(n1255), .A1(n4048), .B0(n3088), .B1(n4060), .Y(n2495) );
  OAI22XL U4012 ( .A0(n1256), .A1(n4048), .B0(n3152), .B1(n4060), .Y(n2496) );
  OAI22XL U4013 ( .A0(n1257), .A1(n4048), .B0(n3151), .B1(n4060), .Y(n2497) );
  OAI22XL U4014 ( .A0(n1258), .A1(n4048), .B0(n3168), .B1(n4060), .Y(n2498) );
  OAI22XL U4015 ( .A0(n1259), .A1(n4048), .B0(n3170), .B1(n4061), .Y(n2499) );
  OAI22XL U4016 ( .A0(n1260), .A1(n4048), .B0(n3159), .B1(n4061), .Y(n2500) );
  OAI22XL U4017 ( .A0(n1261), .A1(n4048), .B0(n3150), .B1(n4061), .Y(n2501) );
  OAI22XL U4018 ( .A0(n1262), .A1(n4048), .B0(n3161), .B1(n4061), .Y(n2502) );
  OAI22XL U4019 ( .A0(n1263), .A1(n4048), .B0(n3149), .B1(n4061), .Y(n2503) );
  OAI22XL U4020 ( .A0(n1264), .A1(n4049), .B0(n3163), .B1(n4061), .Y(n2504) );
  OAI22XL U4021 ( .A0(n1265), .A1(n4049), .B0(n3165), .B1(n4061), .Y(n2505) );
  OAI22XL U4022 ( .A0(n1266), .A1(n4049), .B0(n3167), .B1(n4061), .Y(n2506) );
  OAI22XL U4023 ( .A0(n1267), .A1(n4049), .B0(n3169), .B1(n4061), .Y(n2507) );
  OAI22XL U4024 ( .A0(n1268), .A1(n4049), .B0(n3148), .B1(n4061), .Y(n2508) );
  OAI22XL U4025 ( .A0(n1269), .A1(n4049), .B0(n3147), .B1(n4061), .Y(n2509) );
  OAI22XL U4026 ( .A0(n1270), .A1(n4049), .B0(n3158), .B1(n4062), .Y(n2510) );
  OAI22XL U4027 ( .A0(n1271), .A1(n4049), .B0(n3157), .B1(n4062), .Y(n2511) );
  OAI22XL U4028 ( .A0(n1272), .A1(n4049), .B0(n3166), .B1(n4062), .Y(n2512) );
  OAI22XL U4029 ( .A0(n1273), .A1(n4049), .B0(n3156), .B1(n4062), .Y(n2513) );
  OAI22XL U4030 ( .A0(n1274), .A1(n4049), .B0(n3160), .B1(n4062), .Y(n2514) );
  OAI22XL U4031 ( .A0(n1275), .A1(n4049), .B0(n3162), .B1(n4062), .Y(n2515) );
  OAI22XL U4032 ( .A0(n1276), .A1(n4050), .B0(n3164), .B1(n4062), .Y(n2516) );
  OAI22XL U4033 ( .A0(n1277), .A1(n4050), .B0(n3155), .B1(n4062), .Y(n2517) );
  OAI22XL U4034 ( .A0(n1278), .A1(n4050), .B0(n3154), .B1(n4062), .Y(n2518) );
  OAI22XL U4035 ( .A0(n1279), .A1(n4050), .B0(n3153), .B1(n4062), .Y(n2519) );
  OAI22XL U4036 ( .A0(n1280), .A1(n4050), .B0(n3097), .B1(n4062), .Y(n2520) );
  OAI22XL U4037 ( .A0(n1281), .A1(n4050), .B0(n3093), .B1(n4063), .Y(n2521) );
  OAI22XL U4038 ( .A0(n1282), .A1(n4050), .B0(n3092), .B1(n4063), .Y(n2522) );
  OAI22XL U4039 ( .A0(n1283), .A1(n4050), .B0(n3091), .B1(n4063), .Y(n2523) );
  OAI22XL U4040 ( .A0(n1284), .A1(n4050), .B0(n3090), .B1(n4063), .Y(n2524) );
  OAI22XL U4041 ( .A0(n1285), .A1(n4050), .B0(n3096), .B1(n4063), .Y(n2525) );
  OAI22XL U4042 ( .A0(n1286), .A1(n4050), .B0(n3095), .B1(n4063), .Y(n2526) );
  OAI22XL U4043 ( .A0(n1287), .A1(n4050), .B0(n3094), .B1(n4063), .Y(n2527) );
  OAI22XL U4044 ( .A0(n1288), .A1(n4051), .B0(n3179), .B1(n4063), .Y(n2528) );
  OAI22XL U4045 ( .A0(n1289), .A1(n4051), .B0(n3178), .B1(n4063), .Y(n2529) );
  OAI22XL U4046 ( .A0(n1290), .A1(n4051), .B0(n3177), .B1(n4063), .Y(n2530) );
  OAI22XL U4047 ( .A0(n1291), .A1(n4051), .B0(n3176), .B1(n4063), .Y(n2531) );
  OAI22XL U4048 ( .A0(n1292), .A1(n4051), .B0(n3187), .B1(n4064), .Y(n2532) );
  OAI22XL U4049 ( .A0(n1293), .A1(n4051), .B0(n3186), .B1(n4064), .Y(n2533) );
  OAI22XL U4050 ( .A0(n1294), .A1(n4051), .B0(n3185), .B1(n4064), .Y(n2534) );
  OAI22XL U4051 ( .A0(n1295), .A1(n4051), .B0(n3184), .B1(n4064), .Y(n2535) );
  OAI22XL U4052 ( .A0(n1296), .A1(n4051), .B0(n3183), .B1(n4064), .Y(n2536) );
  OAI22XL U4053 ( .A0(n1297), .A1(n4051), .B0(n3182), .B1(n4064), .Y(n2537) );
  OAI22XL U4054 ( .A0(n1298), .A1(n4051), .B0(n3146), .B1(n4064), .Y(n2538) );
  OAI22XL U4055 ( .A0(n1299), .A1(n4051), .B0(n3145), .B1(n4064), .Y(n2539) );
  OAI22XL U4056 ( .A0(n1300), .A1(n4052), .B0(n3144), .B1(n4064), .Y(n2540) );
  OAI22XL U4057 ( .A0(n1301), .A1(n4052), .B0(n3143), .B1(n4064), .Y(n2541) );
  OAI22XL U4058 ( .A0(n1302), .A1(n4052), .B0(n3142), .B1(n4064), .Y(n2542) );
  OAI22XL U4059 ( .A0(n1303), .A1(n4052), .B0(n3139), .B1(n4065), .Y(n2543) );
  OAI22XL U4060 ( .A0(n1304), .A1(n4052), .B0(n3138), .B1(n4065), .Y(n2544) );
  OAI22XL U4061 ( .A0(n1305), .A1(n4052), .B0(n3137), .B1(n4065), .Y(n2545) );
  OAI22XL U4062 ( .A0(n1306), .A1(n4052), .B0(n3136), .B1(n4065), .Y(n2546) );
  OAI22XL U4063 ( .A0(n1307), .A1(n4052), .B0(n3141), .B1(n4065), .Y(n2547) );
  OAI22XL U4064 ( .A0(n1308), .A1(n4052), .B0(n3135), .B1(n4065), .Y(n2548) );
  OAI22XL U4065 ( .A0(n1309), .A1(n4052), .B0(n3140), .B1(n4065), .Y(n2549) );
  OAI22XL U4066 ( .A0(n1310), .A1(n4052), .B0(n3172), .B1(n4065), .Y(n2550) );
  OAI22XL U4067 ( .A0(n1311), .A1(n4052), .B0(n3180), .B1(n4065), .Y(n2551) );
  OAI22XL U4068 ( .A0(n1312), .A1(n4053), .B0(n3173), .B1(n4065), .Y(n2552) );
  OAI22XL U4069 ( .A0(n1313), .A1(n4053), .B0(n3171), .B1(n4065), .Y(n2553) );
  OAI22XL U4070 ( .A0(n1314), .A1(n4053), .B0(n3189), .B1(n4066), .Y(n2554) );
  OAI22XL U4071 ( .A0(n1315), .A1(n4053), .B0(n3188), .B1(n4066), .Y(n2555) );
  OAI22XL U4072 ( .A0(n1316), .A1(n4053), .B0(n3175), .B1(n4066), .Y(n2556) );
  OAI22XL U4073 ( .A0(n1317), .A1(n4053), .B0(n3181), .B1(n4066), .Y(n2557) );
  OAI22XL U4074 ( .A0(n1318), .A1(n4053), .B0(n3174), .B1(n4066), .Y(n2558) );
  OAI22XL U4075 ( .A0(n1347), .A1(n4015), .B0(n3080), .B1(n4040), .Y(n2587) );
  OAI22XL U4076 ( .A0(n1348), .A1(n4015), .B0(n211), .B1(n4038), .Y(n2588) );
  OAI22XL U4077 ( .A0(n1349), .A1(n4015), .B0(n3081), .B1(n4029), .Y(n2589) );
  OAI22XL U4078 ( .A0(n1350), .A1(n4015), .B0(n3079), .B1(n4039), .Y(n2590) );
  OAI22XL U4079 ( .A0(n1351), .A1(n4015), .B0(n3078), .B1(n4028), .Y(n2591) );
  OAI22XL U4080 ( .A0(n1352), .A1(n4015), .B0(n3077), .B1(n4028), .Y(n2592) );
  OAI22XL U4081 ( .A0(n1353), .A1(n4015), .B0(n3076), .B1(n4028), .Y(n2593) );
  OAI22XL U4082 ( .A0(n1354), .A1(n4015), .B0(n3086), .B1(n4028), .Y(n2594) );
  OAI22XL U4083 ( .A0(n1355), .A1(n4015), .B0(n3085), .B1(n4028), .Y(n2595) );
  OAI22XL U4084 ( .A0(n1356), .A1(n4015), .B0(n3084), .B1(n4028), .Y(n2596) );
  OAI22XL U4085 ( .A0(n1357), .A1(n4015), .B0(n3083), .B1(n4028), .Y(n2597) );
  OAI22XL U4086 ( .A0(n1358), .A1(n4015), .B0(n3082), .B1(n4028), .Y(n2598) );
  OAI22XL U4087 ( .A0(n1359), .A1(n4016), .B0(n222), .B1(n4029), .Y(n2599) );
  OAI22XL U4088 ( .A0(n1360), .A1(n4016), .B0(n223), .B1(n4029), .Y(n2600) );
  OAI22XL U4089 ( .A0(n1361), .A1(n4016), .B0(n3130), .B1(n4029), .Y(n2601) );
  OAI22XL U4090 ( .A0(n1362), .A1(n4016), .B0(n3129), .B1(n4029), .Y(n2602) );
  OAI22XL U4091 ( .A0(n1363), .A1(n4016), .B0(n3128), .B1(n4029), .Y(n2603) );
  OAI22XL U4092 ( .A0(n1364), .A1(n4016), .B0(n3127), .B1(n4029), .Y(n2604) );
  OAI22XL U4093 ( .A0(n1365), .A1(n4016), .B0(n3126), .B1(n4029), .Y(n2605) );
  OAI22XL U4094 ( .A0(n1366), .A1(n4016), .B0(n229), .B1(n4029), .Y(n2606) );
  OAI22XL U4095 ( .A0(n1367), .A1(n4016), .B0(n3134), .B1(n4029), .Y(n2607) );
  OAI22XL U4096 ( .A0(n1368), .A1(n4016), .B0(n3133), .B1(n4029), .Y(n2608) );
  OAI22XL U4097 ( .A0(n1369), .A1(n4016), .B0(n3132), .B1(n4029), .Y(n2609) );
  OAI22XL U4098 ( .A0(n1370), .A1(n4016), .B0(n3131), .B1(n4030), .Y(n2610) );
  OAI22XL U4099 ( .A0(n1371), .A1(n4017), .B0(n3074), .B1(n4030), .Y(n2611) );
  OAI22XL U4100 ( .A0(n1372), .A1(n4017), .B0(n3068), .B1(n4030), .Y(n2612) );
  OAI22XL U4101 ( .A0(n1373), .A1(n4017), .B0(n3065), .B1(n4030), .Y(n2613) );
  OAI22XL U4102 ( .A0(n1374), .A1(n4017), .B0(n3071), .B1(n4030), .Y(n2614) );
  OAI22XL U4103 ( .A0(n1375), .A1(n4017), .B0(n3062), .B1(n4030), .Y(n2615) );
  OAI22XL U4104 ( .A0(n1376), .A1(n4017), .B0(n3059), .B1(n4030), .Y(n2616) );
  OAI22XL U4105 ( .A0(n1377), .A1(n4017), .B0(n3056), .B1(n4030), .Y(n2617) );
  OAI22XL U4106 ( .A0(n1378), .A1(n4017), .B0(n3053), .B1(n4030), .Y(n2618) );
  OAI22XL U4107 ( .A0(n1379), .A1(n4017), .B0(n242), .B1(n4030), .Y(n2619) );
  OAI22XL U4108 ( .A0(n1380), .A1(n4017), .B0(n3125), .B1(n4030), .Y(n2620) );
  OAI22XL U4109 ( .A0(n1381), .A1(n4017), .B0(n3124), .B1(n4031), .Y(n2621) );
  OAI22XL U4110 ( .A0(n1382), .A1(n4017), .B0(n3123), .B1(n4031), .Y(n2622) );
  OAI22XL U4111 ( .A0(n1383), .A1(n4018), .B0(n246), .B1(n4031), .Y(n2623) );
  OAI22XL U4112 ( .A0(n1384), .A1(n4018), .B0(n3122), .B1(n4031), .Y(n2624) );
  OAI22XL U4113 ( .A0(n1385), .A1(n4018), .B0(n3121), .B1(n4031), .Y(n2625) );
  OAI22XL U4114 ( .A0(n1386), .A1(n4018), .B0(n3120), .B1(n4031), .Y(n2626) );
  OAI22XL U4115 ( .A0(n1387), .A1(n4018), .B0(n3119), .B1(n4031), .Y(n2627) );
  OAI22XL U4116 ( .A0(n1388), .A1(n4018), .B0(n3118), .B1(n4031), .Y(n2628) );
  OAI22XL U4117 ( .A0(n1389), .A1(n4018), .B0(n3117), .B1(n4031), .Y(n2629) );
  OAI22XL U4118 ( .A0(n1390), .A1(n4018), .B0(n3116), .B1(n4031), .Y(n2630) );
  OAI22XL U4119 ( .A0(n1391), .A1(n4018), .B0(n3115), .B1(n4031), .Y(n2631) );
  OAI22XL U4120 ( .A0(n1392), .A1(n4018), .B0(n3114), .B1(n4032), .Y(n2632) );
  OAI22XL U4121 ( .A0(n1393), .A1(n4018), .B0(n3113), .B1(n4032), .Y(n2633) );
  OAI22XL U4122 ( .A0(n1394), .A1(n4018), .B0(n3112), .B1(n4032), .Y(n2634) );
  OAI22XL U4123 ( .A0(n1395), .A1(n4019), .B0(n3111), .B1(n4032), .Y(n2635) );
  OAI22XL U4124 ( .A0(n1396), .A1(n4019), .B0(n3110), .B1(n4032), .Y(n2636) );
  OAI22XL U4125 ( .A0(n1397), .A1(n4019), .B0(n3109), .B1(n4032), .Y(n2637) );
  OAI22XL U4126 ( .A0(n1398), .A1(n4019), .B0(n3108), .B1(n4032), .Y(n2638) );
  OAI22XL U4127 ( .A0(n1399), .A1(n4019), .B0(n3107), .B1(n4032), .Y(n2639) );
  OAI22XL U4128 ( .A0(n1400), .A1(n4019), .B0(n3106), .B1(n4032), .Y(n2640) );
  OAI22XL U4129 ( .A0(n1401), .A1(n4019), .B0(n3105), .B1(n4032), .Y(n2641) );
  OAI22XL U4130 ( .A0(n1402), .A1(n4019), .B0(n3104), .B1(n4032), .Y(n2642) );
  OAI22XL U4131 ( .A0(n1403), .A1(n4019), .B0(n3103), .B1(n4033), .Y(n2643) );
  OAI22XL U4132 ( .A0(n1404), .A1(n4019), .B0(n3102), .B1(n4033), .Y(n2644) );
  OAI22XL U4133 ( .A0(n1405), .A1(n4019), .B0(n3089), .B1(n4033), .Y(n2645) );
  OAI22XL U4134 ( .A0(n1406), .A1(n4019), .B0(n3101), .B1(n4033), .Y(n2646) );
  OAI22XL U4135 ( .A0(n1407), .A1(n4020), .B0(n3100), .B1(n4033), .Y(n2647) );
  OAI22XL U4136 ( .A0(n1408), .A1(n4020), .B0(n3099), .B1(n4033), .Y(n2648) );
  OAI22XL U4137 ( .A0(n1409), .A1(n4020), .B0(n3098), .B1(n4033), .Y(n2649) );
  OAI22XL U4138 ( .A0(n1410), .A1(n4020), .B0(n3088), .B1(n4033), .Y(n2650) );
  OAI22XL U4139 ( .A0(n1411), .A1(n4020), .B0(n3152), .B1(n4033), .Y(n2651) );
  OAI22XL U4140 ( .A0(n1412), .A1(n4020), .B0(n3151), .B1(n4033), .Y(n2652) );
  OAI22XL U4141 ( .A0(n1413), .A1(n4020), .B0(n3168), .B1(n4033), .Y(n2653) );
  OAI22XL U4142 ( .A0(n1414), .A1(n4020), .B0(n3170), .B1(n4034), .Y(n2654) );
  OAI22XL U4143 ( .A0(n1415), .A1(n4020), .B0(n3159), .B1(n4034), .Y(n2655) );
  OAI22XL U4144 ( .A0(n1416), .A1(n4020), .B0(n3150), .B1(n4034), .Y(n2656) );
  OAI22XL U4145 ( .A0(n1417), .A1(n4020), .B0(n3161), .B1(n4034), .Y(n2657) );
  OAI22XL U4146 ( .A0(n1418), .A1(n4020), .B0(n3149), .B1(n4034), .Y(n2658) );
  OAI22XL U4147 ( .A0(n1419), .A1(n4021), .B0(n3163), .B1(n4034), .Y(n2659) );
  OAI22XL U4148 ( .A0(n1420), .A1(n4021), .B0(n3165), .B1(n4034), .Y(n2660) );
  OAI22XL U4149 ( .A0(n1421), .A1(n4021), .B0(n3167), .B1(n4034), .Y(n2661) );
  OAI22XL U4150 ( .A0(n1422), .A1(n4021), .B0(n3169), .B1(n4034), .Y(n2662) );
  OAI22XL U4151 ( .A0(n1423), .A1(n4021), .B0(n3148), .B1(n4034), .Y(n2663) );
  OAI22XL U4152 ( .A0(n1424), .A1(n4021), .B0(n3147), .B1(n4034), .Y(n2664) );
  OAI22XL U4153 ( .A0(n1425), .A1(n4021), .B0(n3158), .B1(n4035), .Y(n2665) );
  OAI22XL U4154 ( .A0(n1426), .A1(n4021), .B0(n3157), .B1(n4035), .Y(n2666) );
  OAI22XL U4155 ( .A0(n1427), .A1(n4021), .B0(n3166), .B1(n4035), .Y(n2667) );
  OAI22XL U4156 ( .A0(n1428), .A1(n4021), .B0(n3156), .B1(n4035), .Y(n2668) );
  OAI22XL U4157 ( .A0(n1429), .A1(n4021), .B0(n3160), .B1(n4035), .Y(n2669) );
  OAI22XL U4158 ( .A0(n1430), .A1(n4021), .B0(n3162), .B1(n4035), .Y(n2670) );
  OAI22XL U4159 ( .A0(n1431), .A1(n4022), .B0(n3164), .B1(n4035), .Y(n2671) );
  OAI22XL U4160 ( .A0(n1432), .A1(n4022), .B0(n3155), .B1(n4035), .Y(n2672) );
  OAI22XL U4161 ( .A0(n1433), .A1(n4022), .B0(n3154), .B1(n4035), .Y(n2673) );
  OAI22XL U4162 ( .A0(n1434), .A1(n4022), .B0(n3153), .B1(n4035), .Y(n2674) );
  OAI22XL U4163 ( .A0(n1435), .A1(n4022), .B0(n3097), .B1(n4035), .Y(n2675) );
  OAI22XL U4164 ( .A0(n1436), .A1(n4022), .B0(n3093), .B1(n4036), .Y(n2676) );
  OAI22XL U4165 ( .A0(n1437), .A1(n4022), .B0(n3092), .B1(n4036), .Y(n2677) );
  OAI22XL U4166 ( .A0(n1438), .A1(n4022), .B0(n3091), .B1(n4036), .Y(n2678) );
  OAI22XL U4167 ( .A0(n1439), .A1(n4022), .B0(n3090), .B1(n4036), .Y(n2679) );
  OAI22XL U4168 ( .A0(n1440), .A1(n4022), .B0(n3096), .B1(n4036), .Y(n2680) );
  OAI22XL U4169 ( .A0(n1441), .A1(n4022), .B0(n3095), .B1(n4036), .Y(n2681) );
  OAI22XL U4170 ( .A0(n1442), .A1(n4022), .B0(n3094), .B1(n4036), .Y(n2682) );
  OAI22XL U4171 ( .A0(n1443), .A1(n4023), .B0(n3179), .B1(n4036), .Y(n2683) );
  OAI22XL U4172 ( .A0(n1444), .A1(n4023), .B0(n3178), .B1(n4036), .Y(n2684) );
  OAI22XL U4173 ( .A0(n1445), .A1(n4023), .B0(n3177), .B1(n4036), .Y(n2685) );
  OAI22XL U4174 ( .A0(n1446), .A1(n4023), .B0(n3176), .B1(n4036), .Y(n2686) );
  OAI22XL U4175 ( .A0(n1447), .A1(n4023), .B0(n3187), .B1(n4037), .Y(n2687) );
  OAI22XL U4176 ( .A0(n1448), .A1(n4023), .B0(n3186), .B1(n4037), .Y(n2688) );
  OAI22XL U4177 ( .A0(n1449), .A1(n4023), .B0(n3185), .B1(n4037), .Y(n2689) );
  OAI22XL U4178 ( .A0(n1450), .A1(n4023), .B0(n3184), .B1(n4037), .Y(n2690) );
  OAI22XL U4179 ( .A0(n1451), .A1(n4023), .B0(n3183), .B1(n4037), .Y(n2691) );
  OAI22XL U4180 ( .A0(n1452), .A1(n4023), .B0(n3182), .B1(n4037), .Y(n2692) );
  OAI22XL U4181 ( .A0(n1453), .A1(n4023), .B0(n3146), .B1(n4037), .Y(n2693) );
  OAI22XL U4182 ( .A0(n1454), .A1(n4023), .B0(n3145), .B1(n4037), .Y(n2694) );
  OAI22XL U4183 ( .A0(n1455), .A1(n4024), .B0(n3144), .B1(n4037), .Y(n2695) );
  OAI22XL U4184 ( .A0(n1456), .A1(n4024), .B0(n3143), .B1(n4037), .Y(n2696) );
  OAI22XL U4185 ( .A0(n1457), .A1(n4024), .B0(n3142), .B1(n4037), .Y(n2697) );
  OAI22XL U4186 ( .A0(n1458), .A1(n4024), .B0(n3139), .B1(n4038), .Y(n2698) );
  OAI22XL U4187 ( .A0(n1459), .A1(n4024), .B0(n3138), .B1(n4038), .Y(n2699) );
  OAI22XL U4188 ( .A0(n1460), .A1(n4024), .B0(n3137), .B1(n4038), .Y(n2700) );
  OAI22XL U4189 ( .A0(n1461), .A1(n4024), .B0(n3136), .B1(n4038), .Y(n2701) );
  OAI22XL U4190 ( .A0(n1462), .A1(n4024), .B0(n3141), .B1(n4038), .Y(n2702) );
  OAI22XL U4191 ( .A0(n1463), .A1(n4024), .B0(n3135), .B1(n4038), .Y(n2703) );
  OAI22XL U4192 ( .A0(n1464), .A1(n4024), .B0(n3140), .B1(n4038), .Y(n2704) );
  OAI22XL U4193 ( .A0(n1465), .A1(n4024), .B0(n3172), .B1(n4038), .Y(n2705) );
  OAI22XL U4194 ( .A0(n1466), .A1(n4024), .B0(n3180), .B1(n4038), .Y(n2706) );
  OAI22XL U4195 ( .A0(n1467), .A1(n4025), .B0(n3173), .B1(n4038), .Y(n2707) );
  OAI22XL U4196 ( .A0(n1468), .A1(n4025), .B0(n3171), .B1(n4038), .Y(n2708) );
  OAI22XL U4197 ( .A0(n1469), .A1(n4025), .B0(n3189), .B1(n4029), .Y(n2709) );
  OAI22XL U4198 ( .A0(n1470), .A1(n4025), .B0(n3188), .B1(n4040), .Y(n2710) );
  OAI22XL U4199 ( .A0(n1471), .A1(n4025), .B0(n3175), .B1(n4030), .Y(n2711) );
  OAI22XL U4200 ( .A0(n1472), .A1(n4025), .B0(n3181), .B1(n4031), .Y(n2712) );
  OAI22XL U4201 ( .A0(n1473), .A1(n4025), .B0(n3174), .B1(n4034), .Y(n2713) );
  OAI22XL U4202 ( .A0(n1502), .A1(n3987), .B0(n3080), .B1(n4012), .Y(n2742) );
  OAI22XL U4203 ( .A0(n1503), .A1(n3987), .B0(n211), .B1(n3999), .Y(n2743) );
  OAI22XL U4204 ( .A0(n1504), .A1(n3987), .B0(n3081), .B1(n4009), .Y(n2744) );
  OAI22XL U4205 ( .A0(n1505), .A1(n3987), .B0(n3079), .B1(n4011), .Y(n2745) );
  OAI22XL U4206 ( .A0(n1506), .A1(n3987), .B0(n3078), .B1(n4004), .Y(n2746) );
  OAI22XL U4207 ( .A0(n1507), .A1(n3987), .B0(n3077), .B1(n4007), .Y(n2747) );
  OAI22XL U4208 ( .A0(n1508), .A1(n3987), .B0(n3076), .B1(n4003), .Y(n2748) );
  OAI22XL U4209 ( .A0(n1509), .A1(n3987), .B0(n3086), .B1(n4004), .Y(n2749) );
  OAI22XL U4210 ( .A0(n1510), .A1(n3987), .B0(n3085), .B1(n4007), .Y(n2750) );
  OAI22XL U4211 ( .A0(n1511), .A1(n3987), .B0(n3084), .B1(n4003), .Y(n2751) );
  OAI22XL U4212 ( .A0(n1512), .A1(n3987), .B0(n3083), .B1(n4011), .Y(n2752) );
  OAI22XL U4213 ( .A0(n1513), .A1(n3987), .B0(n3082), .B1(n4012), .Y(n2753) );
  OAI22XL U4214 ( .A0(n1514), .A1(n3988), .B0(n222), .B1(n4000), .Y(n2754) );
  OAI22XL U4215 ( .A0(n1515), .A1(n3988), .B0(n223), .B1(n4000), .Y(n2755) );
  OAI22XL U4216 ( .A0(n1516), .A1(n3988), .B0(n3130), .B1(n4000), .Y(n2756) );
  OAI22XL U4217 ( .A0(n1517), .A1(n3988), .B0(n3129), .B1(n4000), .Y(n2757) );
  OAI22XL U4218 ( .A0(n1518), .A1(n3988), .B0(n3128), .B1(n4000), .Y(n2758) );
  OAI22XL U4219 ( .A0(n1519), .A1(n3988), .B0(n3127), .B1(n4000), .Y(n2759) );
  OAI22XL U4220 ( .A0(n1520), .A1(n3988), .B0(n3126), .B1(n4000), .Y(n2760) );
  OAI22XL U4221 ( .A0(n1521), .A1(n3988), .B0(n229), .B1(n4000), .Y(n2761) );
  OAI22XL U4222 ( .A0(n1522), .A1(n3988), .B0(n3134), .B1(n4000), .Y(n2762) );
  OAI22XL U4223 ( .A0(n1523), .A1(n3988), .B0(n3133), .B1(n4000), .Y(n2763) );
  OAI22XL U4224 ( .A0(n1524), .A1(n3988), .B0(n3132), .B1(n4000), .Y(n2764) );
  OAI22XL U4225 ( .A0(n1525), .A1(n3988), .B0(n3131), .B1(n4001), .Y(n2765) );
  OAI22XL U4226 ( .A0(n1526), .A1(n3989), .B0(n3073), .B1(n4001), .Y(n2766) );
  OAI22XL U4227 ( .A0(n1527), .A1(n3989), .B0(n3067), .B1(n4001), .Y(n2767) );
  OAI22XL U4228 ( .A0(n1528), .A1(n3989), .B0(n3064), .B1(n4001), .Y(n2768) );
  OAI22XL U4229 ( .A0(n1529), .A1(n3989), .B0(n3070), .B1(n4001), .Y(n2769) );
  OAI22XL U4230 ( .A0(n1530), .A1(n3989), .B0(n3061), .B1(n4001), .Y(n2770) );
  OAI22XL U4231 ( .A0(n1531), .A1(n3989), .B0(n3058), .B1(n4001), .Y(n2771) );
  OAI22XL U4232 ( .A0(n1532), .A1(n3989), .B0(n3055), .B1(n4001), .Y(n2772) );
  OAI22XL U4233 ( .A0(n1533), .A1(n3989), .B0(n3053), .B1(n4001), .Y(n2773) );
  OAI22XL U4234 ( .A0(n1534), .A1(n3989), .B0(n242), .B1(n4001), .Y(n2774) );
  OAI22XL U4235 ( .A0(n1535), .A1(n3989), .B0(n3125), .B1(n4001), .Y(n2775) );
  OAI22XL U4236 ( .A0(n1536), .A1(n3989), .B0(n3124), .B1(n4002), .Y(n2776) );
  OAI22XL U4237 ( .A0(n1537), .A1(n3989), .B0(n3123), .B1(n4002), .Y(n2777) );
  OAI22XL U4238 ( .A0(n1538), .A1(n3990), .B0(n246), .B1(n4002), .Y(n2778) );
  OAI22XL U4239 ( .A0(n1539), .A1(n3990), .B0(n3122), .B1(n4002), .Y(n2779) );
  OAI22XL U4240 ( .A0(n1540), .A1(n3990), .B0(n3121), .B1(n4002), .Y(n2780) );
  OAI22XL U4241 ( .A0(n1541), .A1(n3990), .B0(n3120), .B1(n4002), .Y(n2781) );
  OAI22XL U4242 ( .A0(n1542), .A1(n3990), .B0(n3119), .B1(n4002), .Y(n2782) );
  OAI22XL U4243 ( .A0(n1543), .A1(n3990), .B0(n3118), .B1(n4002), .Y(n2783) );
  OAI22XL U4244 ( .A0(n1544), .A1(n3990), .B0(n3117), .B1(n4002), .Y(n2784) );
  OAI22XL U4245 ( .A0(n1545), .A1(n3990), .B0(n3116), .B1(n4002), .Y(n2785) );
  OAI22XL U4246 ( .A0(n1546), .A1(n3990), .B0(n3115), .B1(n4002), .Y(n2786) );
  OAI22XL U4247 ( .A0(n1547), .A1(n3990), .B0(n3114), .B1(n4003), .Y(n2787) );
  OAI22XL U4248 ( .A0(n1548), .A1(n3990), .B0(n3113), .B1(n4003), .Y(n2788) );
  OAI22XL U4249 ( .A0(n1549), .A1(n3990), .B0(n3112), .B1(n4003), .Y(n2789) );
  OAI22XL U4250 ( .A0(n1550), .A1(n3991), .B0(n3111), .B1(n4003), .Y(n2790) );
  OAI22XL U4251 ( .A0(n1551), .A1(n3991), .B0(n3110), .B1(n4003), .Y(n2791) );
  OAI22XL U4252 ( .A0(n1552), .A1(n3991), .B0(n3109), .B1(n4003), .Y(n2792) );
  OAI22XL U4253 ( .A0(n1553), .A1(n3991), .B0(n3108), .B1(n4003), .Y(n2793) );
  OAI22XL U4254 ( .A0(n1554), .A1(n3991), .B0(n3107), .B1(n4003), .Y(n2794) );
  OAI22XL U4255 ( .A0(n1555), .A1(n3991), .B0(n3106), .B1(n4003), .Y(n2795) );
  OAI22XL U4256 ( .A0(n1556), .A1(n3991), .B0(n3105), .B1(n4003), .Y(n2796) );
  OAI22XL U4257 ( .A0(n1557), .A1(n3991), .B0(n3104), .B1(n4003), .Y(n2797) );
  OAI22XL U4258 ( .A0(n1558), .A1(n3991), .B0(n3103), .B1(n4004), .Y(n2798) );
  OAI22XL U4259 ( .A0(n1559), .A1(n3991), .B0(n3102), .B1(n4004), .Y(n2799) );
  OAI22XL U4260 ( .A0(n1560), .A1(n3991), .B0(n3089), .B1(n4004), .Y(n2800) );
  OAI22XL U4261 ( .A0(n1561), .A1(n3991), .B0(n3101), .B1(n4004), .Y(n2801) );
  OAI22XL U4262 ( .A0(n1562), .A1(n3992), .B0(n3100), .B1(n4004), .Y(n2802) );
  OAI22XL U4263 ( .A0(n1563), .A1(n3992), .B0(n3099), .B1(n4004), .Y(n2803) );
  OAI22XL U4264 ( .A0(n1564), .A1(n3992), .B0(n3098), .B1(n4004), .Y(n2804) );
  OAI22XL U4265 ( .A0(n1565), .A1(n3992), .B0(n3088), .B1(n4004), .Y(n2805) );
  OAI22XL U4266 ( .A0(n1566), .A1(n3992), .B0(n3152), .B1(n4004), .Y(n2806) );
  OAI22XL U4267 ( .A0(n1567), .A1(n3992), .B0(n3151), .B1(n4004), .Y(n2807) );
  OAI22XL U4268 ( .A0(n1568), .A1(n3992), .B0(n3168), .B1(n4004), .Y(n2808) );
  OAI22XL U4269 ( .A0(n1569), .A1(n3992), .B0(n3170), .B1(n4005), .Y(n2809) );
  OAI22XL U4270 ( .A0(n1570), .A1(n3992), .B0(n3159), .B1(n4005), .Y(n2810) );
  OAI22XL U4271 ( .A0(n1571), .A1(n3992), .B0(n3150), .B1(n4005), .Y(n2811) );
  OAI22XL U4272 ( .A0(n1572), .A1(n3992), .B0(n3161), .B1(n4005), .Y(n2812) );
  OAI22XL U4273 ( .A0(n1573), .A1(n3992), .B0(n3149), .B1(n4005), .Y(n2813) );
  OAI22XL U4274 ( .A0(n1574), .A1(n3993), .B0(n3163), .B1(n4005), .Y(n2814) );
  OAI22XL U4275 ( .A0(n1575), .A1(n3993), .B0(n3165), .B1(n4005), .Y(n2815) );
  OAI22XL U4276 ( .A0(n1576), .A1(n3993), .B0(n3167), .B1(n4005), .Y(n2816) );
  OAI22XL U4277 ( .A0(n1577), .A1(n3993), .B0(n3169), .B1(n4005), .Y(n2817) );
  OAI22XL U4278 ( .A0(n1578), .A1(n3993), .B0(n3148), .B1(n4005), .Y(n2818) );
  OAI22XL U4279 ( .A0(n1579), .A1(n3993), .B0(n3147), .B1(n4005), .Y(n2819) );
  OAI22XL U4280 ( .A0(n1580), .A1(n3993), .B0(n3158), .B1(n4006), .Y(n2820) );
  OAI22XL U4281 ( .A0(n1581), .A1(n3993), .B0(n3157), .B1(n4006), .Y(n2821) );
  OAI22XL U4282 ( .A0(n1582), .A1(n3993), .B0(n3166), .B1(n4006), .Y(n2822) );
  OAI22XL U4283 ( .A0(n1583), .A1(n3993), .B0(n3156), .B1(n4006), .Y(n2823) );
  OAI22XL U4284 ( .A0(n1584), .A1(n3993), .B0(n3160), .B1(n4006), .Y(n2824) );
  OAI22XL U4285 ( .A0(n1585), .A1(n3993), .B0(n3162), .B1(n4006), .Y(n2825) );
  OAI22XL U4286 ( .A0(n1586), .A1(n3994), .B0(n3164), .B1(n4006), .Y(n2826) );
  OAI22XL U4287 ( .A0(n1587), .A1(n3994), .B0(n3155), .B1(n4006), .Y(n2827) );
  OAI22XL U4288 ( .A0(n1588), .A1(n3994), .B0(n3154), .B1(n4006), .Y(n2828) );
  OAI22XL U4289 ( .A0(n1589), .A1(n3994), .B0(n3153), .B1(n4006), .Y(n2829) );
  OAI22XL U4290 ( .A0(n1590), .A1(n3994), .B0(n3097), .B1(n4006), .Y(n2830) );
  OAI22XL U4291 ( .A0(n1591), .A1(n3994), .B0(n3093), .B1(n4007), .Y(n2831) );
  OAI22XL U4292 ( .A0(n1592), .A1(n3994), .B0(n3092), .B1(n4007), .Y(n2832) );
  OAI22XL U4293 ( .A0(n1593), .A1(n3994), .B0(n3091), .B1(n4007), .Y(n2833) );
  OAI22XL U4294 ( .A0(n1594), .A1(n3994), .B0(n3090), .B1(n4007), .Y(n2834) );
  OAI22XL U4295 ( .A0(n1595), .A1(n3994), .B0(n3096), .B1(n4007), .Y(n2835) );
  OAI22XL U4296 ( .A0(n1596), .A1(n3994), .B0(n3095), .B1(n4007), .Y(n2836) );
  OAI22XL U4297 ( .A0(n1597), .A1(n3994), .B0(n3094), .B1(n4007), .Y(n2837) );
  OAI22XL U4298 ( .A0(n1598), .A1(n3995), .B0(n3179), .B1(n4007), .Y(n2838) );
  OAI22XL U4299 ( .A0(n1599), .A1(n3995), .B0(n3178), .B1(n4007), .Y(n2839) );
  OAI22XL U4300 ( .A0(n1600), .A1(n3995), .B0(n3177), .B1(n4007), .Y(n2840) );
  OAI22XL U4301 ( .A0(n1601), .A1(n3995), .B0(n3176), .B1(n4007), .Y(n2841) );
  OAI22XL U4302 ( .A0(n1602), .A1(n3995), .B0(n3187), .B1(n4008), .Y(n2842) );
  OAI22XL U4303 ( .A0(n1603), .A1(n3995), .B0(n3186), .B1(n4008), .Y(n2843) );
  OAI22XL U4304 ( .A0(n1604), .A1(n3995), .B0(n3185), .B1(n4008), .Y(n2844) );
  OAI22XL U4305 ( .A0(n1605), .A1(n3995), .B0(n3184), .B1(n4008), .Y(n2845) );
  OAI22XL U4306 ( .A0(n1606), .A1(n3995), .B0(n3183), .B1(n4008), .Y(n2846) );
  OAI22XL U4307 ( .A0(n1607), .A1(n3995), .B0(n3182), .B1(n4008), .Y(n2847) );
  OAI22XL U4308 ( .A0(n1608), .A1(n3995), .B0(n3146), .B1(n4008), .Y(n2848) );
  OAI22XL U4309 ( .A0(n1609), .A1(n3995), .B0(n3145), .B1(n4008), .Y(n2849) );
  OAI22XL U4310 ( .A0(n1610), .A1(n3996), .B0(n3144), .B1(n4008), .Y(n2850) );
  OAI22XL U4311 ( .A0(n1611), .A1(n3996), .B0(n3143), .B1(n4008), .Y(n2851) );
  OAI22XL U4312 ( .A0(n1612), .A1(n3996), .B0(n3142), .B1(n4008), .Y(n2852) );
  OAI22XL U4313 ( .A0(n1613), .A1(n3996), .B0(n3139), .B1(n4009), .Y(n2853) );
  OAI22XL U4314 ( .A0(n1614), .A1(n3996), .B0(n3138), .B1(n4009), .Y(n2854) );
  OAI22XL U4315 ( .A0(n1615), .A1(n3996), .B0(n3137), .B1(n4009), .Y(n2855) );
  OAI22XL U4316 ( .A0(n1616), .A1(n3996), .B0(n3136), .B1(n4009), .Y(n2856) );
  OAI22XL U4317 ( .A0(n1617), .A1(n3996), .B0(n3141), .B1(n4009), .Y(n2857) );
  OAI22XL U4318 ( .A0(n1618), .A1(n3996), .B0(n3135), .B1(n4009), .Y(n2858) );
  OAI22XL U4319 ( .A0(n1619), .A1(n3996), .B0(n3140), .B1(n4009), .Y(n2859) );
  OAI22XL U4320 ( .A0(n1620), .A1(n3996), .B0(n3172), .B1(n4009), .Y(n2860) );
  OAI22XL U4321 ( .A0(n1621), .A1(n3996), .B0(n3180), .B1(n4009), .Y(n2861) );
  OAI22XL U4322 ( .A0(n1622), .A1(n3997), .B0(n3173), .B1(n4009), .Y(n2862) );
  OAI22XL U4323 ( .A0(n1623), .A1(n3997), .B0(n3171), .B1(n4009), .Y(n2863) );
  OAI22XL U4324 ( .A0(n1624), .A1(n3997), .B0(n3189), .B1(n4010), .Y(n2864) );
  OAI22XL U4325 ( .A0(n1625), .A1(n3997), .B0(n3188), .B1(n4010), .Y(n2865) );
  OAI22XL U4326 ( .A0(n1626), .A1(n3997), .B0(n3175), .B1(n4010), .Y(n2866) );
  OAI22XL U4327 ( .A0(n1627), .A1(n3997), .B0(n3181), .B1(n4010), .Y(n2867) );
  OAI22XL U4328 ( .A0(n1628), .A1(n3997), .B0(n3174), .B1(n4010), .Y(n2868) );
  OAI22XL U4329 ( .A0(n1657), .A1(n3959), .B0(n3080), .B1(n3984), .Y(n2897) );
  OAI22XL U4330 ( .A0(n1658), .A1(n3959), .B0(n211), .B1(n3982), .Y(n2898) );
  OAI22XL U4331 ( .A0(n1659), .A1(n3959), .B0(n3081), .B1(n3973), .Y(n2899) );
  OAI22XL U4332 ( .A0(n1660), .A1(n3959), .B0(n3079), .B1(n3983), .Y(n2900) );
  OAI22XL U4333 ( .A0(n1661), .A1(n3959), .B0(n3078), .B1(n3972), .Y(n2901) );
  OAI22XL U4334 ( .A0(n1662), .A1(n3959), .B0(n3077), .B1(n3972), .Y(n2902) );
  OAI22XL U4335 ( .A0(n1663), .A1(n3959), .B0(n3076), .B1(n3972), .Y(n2903) );
  OAI22XL U4336 ( .A0(n1664), .A1(n3959), .B0(n3086), .B1(n3972), .Y(n2904) );
  OAI22XL U4337 ( .A0(n1665), .A1(n3959), .B0(n3085), .B1(n3972), .Y(n2905) );
  OAI22XL U4338 ( .A0(n1666), .A1(n3959), .B0(n3084), .B1(n3972), .Y(n2906) );
  OAI22XL U4339 ( .A0(n1667), .A1(n3959), .B0(n3083), .B1(n3972), .Y(n2907) );
  OAI22XL U4340 ( .A0(n1668), .A1(n3959), .B0(n3082), .B1(n3972), .Y(n2908) );
  OAI22XL U4341 ( .A0(n1669), .A1(n3960), .B0(n222), .B1(n3973), .Y(n2909) );
  OAI22XL U4342 ( .A0(n1670), .A1(n3960), .B0(n223), .B1(n3973), .Y(n2910) );
  OAI22XL U4343 ( .A0(n1671), .A1(n3960), .B0(n3130), .B1(n3973), .Y(n2911) );
  OAI22XL U4344 ( .A0(n1672), .A1(n3960), .B0(n3129), .B1(n3973), .Y(n2912) );
  OAI22XL U4345 ( .A0(n1673), .A1(n3960), .B0(n3128), .B1(n3973), .Y(n2913) );
  OAI22XL U4346 ( .A0(n1674), .A1(n3960), .B0(n3127), .B1(n3973), .Y(n2914) );
  OAI22XL U4347 ( .A0(n1675), .A1(n3960), .B0(n3126), .B1(n3973), .Y(n2915) );
  OAI22XL U4348 ( .A0(n1676), .A1(n3960), .B0(n229), .B1(n3973), .Y(n2916) );
  OAI22XL U4349 ( .A0(n1677), .A1(n3960), .B0(n3134), .B1(n3973), .Y(n2917) );
  OAI22XL U4350 ( .A0(n1678), .A1(n3960), .B0(n3133), .B1(n3973), .Y(n2918) );
  OAI22XL U4351 ( .A0(n1679), .A1(n3960), .B0(n3132), .B1(n3973), .Y(n2919) );
  OAI22XL U4352 ( .A0(n1680), .A1(n3960), .B0(n3131), .B1(n3974), .Y(n2920) );
  OAI22XL U4353 ( .A0(n1681), .A1(n3961), .B0(n3074), .B1(n3974), .Y(n2921) );
  OAI22XL U4354 ( .A0(n1682), .A1(n3961), .B0(n3068), .B1(n3974), .Y(n2922) );
  OAI22XL U4355 ( .A0(n1683), .A1(n3961), .B0(n3065), .B1(n3974), .Y(n2923) );
  OAI22XL U4356 ( .A0(n1684), .A1(n3961), .B0(n3071), .B1(n3974), .Y(n2924) );
  OAI22XL U4357 ( .A0(n1685), .A1(n3961), .B0(n3062), .B1(n3974), .Y(n2925) );
  OAI22XL U4358 ( .A0(n1686), .A1(n3961), .B0(n3059), .B1(n3974), .Y(n2926) );
  OAI22XL U4359 ( .A0(n1687), .A1(n3961), .B0(n3056), .B1(n3974), .Y(n2927) );
  OAI22XL U4360 ( .A0(n1688), .A1(n3961), .B0(n3053), .B1(n3974), .Y(n2928) );
  OAI22XL U4361 ( .A0(n1689), .A1(n3961), .B0(n242), .B1(n3974), .Y(n2929) );
  OAI22XL U4362 ( .A0(n1690), .A1(n3961), .B0(n3125), .B1(n3974), .Y(n2930) );
  OAI22XL U4363 ( .A0(n1691), .A1(n3961), .B0(n3124), .B1(n3975), .Y(n2931) );
  OAI22XL U4364 ( .A0(n1692), .A1(n3961), .B0(n3123), .B1(n3975), .Y(n2932) );
  OAI22XL U4365 ( .A0(n1693), .A1(n3962), .B0(n246), .B1(n3975), .Y(n2933) );
  OAI22XL U4366 ( .A0(n1694), .A1(n3962), .B0(n3122), .B1(n3975), .Y(n2934) );
  OAI22XL U4367 ( .A0(n1695), .A1(n3962), .B0(n3121), .B1(n3975), .Y(n2935) );
  OAI22XL U4368 ( .A0(n1696), .A1(n3962), .B0(n3120), .B1(n3975), .Y(n2936) );
  OAI22XL U4369 ( .A0(n1697), .A1(n3962), .B0(n3119), .B1(n3975), .Y(n2937) );
  OAI22XL U4370 ( .A0(n1698), .A1(n3962), .B0(n3118), .B1(n3975), .Y(n2938) );
  OAI22XL U4371 ( .A0(n1699), .A1(n3962), .B0(n3117), .B1(n3975), .Y(n2939) );
  OAI22XL U4372 ( .A0(n1700), .A1(n3962), .B0(n3116), .B1(n3975), .Y(n2940) );
  OAI22XL U4373 ( .A0(n1701), .A1(n3962), .B0(n3115), .B1(n3975), .Y(n2941) );
  OAI22XL U4374 ( .A0(n1702), .A1(n3962), .B0(n3114), .B1(n3976), .Y(n2942) );
  OAI22XL U4375 ( .A0(n1703), .A1(n3962), .B0(n3113), .B1(n3976), .Y(n2943) );
  OAI22XL U4376 ( .A0(n1704), .A1(n3962), .B0(n3112), .B1(n3976), .Y(n2944) );
  OAI22XL U4377 ( .A0(n1705), .A1(n3963), .B0(n3111), .B1(n3976), .Y(n2945) );
  OAI22XL U4378 ( .A0(n1706), .A1(n3963), .B0(n3110), .B1(n3976), .Y(n2946) );
  OAI22XL U4379 ( .A0(n1707), .A1(n3963), .B0(n3109), .B1(n3976), .Y(n2947) );
  OAI22XL U4380 ( .A0(n1708), .A1(n3963), .B0(n3108), .B1(n3976), .Y(n2948) );
  OAI22XL U4381 ( .A0(n1709), .A1(n3963), .B0(n3107), .B1(n3976), .Y(n2949) );
  OAI22XL U4382 ( .A0(n1710), .A1(n3963), .B0(n3106), .B1(n3976), .Y(n2950) );
  OAI22XL U4383 ( .A0(n1711), .A1(n3963), .B0(n3105), .B1(n3976), .Y(n2951) );
  OAI22XL U4384 ( .A0(n1712), .A1(n3963), .B0(n3104), .B1(n3976), .Y(n2952) );
  OAI22XL U4385 ( .A0(n1713), .A1(n3963), .B0(n3103), .B1(n3977), .Y(n2953) );
  OAI22XL U4386 ( .A0(n1714), .A1(n3963), .B0(n3102), .B1(n3977), .Y(n2954) );
  OAI22XL U4387 ( .A0(n1715), .A1(n3963), .B0(n3089), .B1(n3977), .Y(n2955) );
  OAI22XL U4388 ( .A0(n1716), .A1(n3963), .B0(n3101), .B1(n3977), .Y(n2956) );
  OAI22XL U4389 ( .A0(n1717), .A1(n3964), .B0(n3100), .B1(n3977), .Y(n2957) );
  OAI22XL U4390 ( .A0(n1718), .A1(n3964), .B0(n3099), .B1(n3977), .Y(n2958) );
  OAI22XL U4391 ( .A0(n1719), .A1(n3964), .B0(n3098), .B1(n3977), .Y(n2959) );
  OAI22XL U4392 ( .A0(n1720), .A1(n3964), .B0(n3088), .B1(n3977), .Y(n2960) );
  OAI22XL U4393 ( .A0(n1721), .A1(n3964), .B0(n3152), .B1(n3977), .Y(n2961) );
  OAI22XL U4394 ( .A0(n1722), .A1(n3964), .B0(n3151), .B1(n3977), .Y(n2962) );
  OAI22XL U4395 ( .A0(n1723), .A1(n3964), .B0(n3168), .B1(n3977), .Y(n2963) );
  OAI22XL U4396 ( .A0(n1724), .A1(n3964), .B0(n3170), .B1(n3978), .Y(n2964) );
  OAI22XL U4397 ( .A0(n1725), .A1(n3964), .B0(n3159), .B1(n3978), .Y(n2965) );
  OAI22XL U4398 ( .A0(n1726), .A1(n3964), .B0(n3150), .B1(n3978), .Y(n2966) );
  OAI22XL U4399 ( .A0(n1727), .A1(n3964), .B0(n3161), .B1(n3978), .Y(n2967) );
  OAI22XL U4400 ( .A0(n1728), .A1(n3964), .B0(n3149), .B1(n3978), .Y(n2968) );
  OAI22XL U4401 ( .A0(n1729), .A1(n3965), .B0(n3163), .B1(n3978), .Y(n2969) );
  OAI22XL U4402 ( .A0(n1730), .A1(n3965), .B0(n3165), .B1(n3978), .Y(n2970) );
  OAI22XL U4403 ( .A0(n1731), .A1(n3965), .B0(n3167), .B1(n3978), .Y(n2971) );
  OAI22XL U4404 ( .A0(n1732), .A1(n3965), .B0(n3169), .B1(n3978), .Y(n2972) );
  OAI22XL U4405 ( .A0(n1733), .A1(n3965), .B0(n3148), .B1(n3978), .Y(n2973) );
  OAI22XL U4406 ( .A0(n1734), .A1(n3965), .B0(n3147), .B1(n3978), .Y(n2974) );
  OAI22XL U4407 ( .A0(n1735), .A1(n3965), .B0(n3158), .B1(n3979), .Y(n2975) );
  OAI22XL U4408 ( .A0(n1736), .A1(n3965), .B0(n3157), .B1(n3979), .Y(n2976) );
  OAI22XL U4409 ( .A0(n1737), .A1(n3965), .B0(n3166), .B1(n3979), .Y(n2977) );
  OAI22XL U4410 ( .A0(n1738), .A1(n3965), .B0(n3156), .B1(n3979), .Y(n2978) );
  OAI22XL U4411 ( .A0(n1739), .A1(n3965), .B0(n3160), .B1(n3979), .Y(n2979) );
  OAI22XL U4412 ( .A0(n1740), .A1(n3965), .B0(n3162), .B1(n3979), .Y(n2980) );
  OAI22XL U4413 ( .A0(n1741), .A1(n3966), .B0(n3164), .B1(n3979), .Y(n2981) );
  OAI22XL U4414 ( .A0(n1742), .A1(n3966), .B0(n3155), .B1(n3979), .Y(n2982) );
  OAI22XL U4415 ( .A0(n1743), .A1(n3966), .B0(n3154), .B1(n3979), .Y(n2983) );
  OAI22XL U4416 ( .A0(n1744), .A1(n3966), .B0(n3153), .B1(n3979), .Y(n2984) );
  OAI22XL U4417 ( .A0(n1745), .A1(n3966), .B0(n3097), .B1(n3979), .Y(n2985) );
  OAI22XL U4418 ( .A0(n1746), .A1(n3966), .B0(n3093), .B1(n3980), .Y(n2986) );
  OAI22XL U4419 ( .A0(n1747), .A1(n3966), .B0(n3092), .B1(n3980), .Y(n2987) );
  OAI22XL U4420 ( .A0(n1748), .A1(n3966), .B0(n3091), .B1(n3980), .Y(n2988) );
  OAI22XL U4421 ( .A0(n1749), .A1(n3966), .B0(n3090), .B1(n3980), .Y(n2989) );
  OAI22XL U4422 ( .A0(n1750), .A1(n3966), .B0(n3096), .B1(n3980), .Y(n2990) );
  OAI22XL U4423 ( .A0(n1751), .A1(n3966), .B0(n3095), .B1(n3980), .Y(n2991) );
  OAI22XL U4424 ( .A0(n1752), .A1(n3966), .B0(n3094), .B1(n3980), .Y(n2992) );
  OAI22XL U4425 ( .A0(n1753), .A1(n3967), .B0(n3179), .B1(n3980), .Y(n2993) );
  OAI22XL U4426 ( .A0(n1754), .A1(n3967), .B0(n3178), .B1(n3980), .Y(n2994) );
  OAI22XL U4427 ( .A0(n1755), .A1(n3967), .B0(n3177), .B1(n3980), .Y(n2995) );
  OAI22XL U4428 ( .A0(n1756), .A1(n3967), .B0(n3176), .B1(n3980), .Y(n2996) );
  OAI22XL U4429 ( .A0(n1757), .A1(n3967), .B0(n3187), .B1(n3981), .Y(n2997) );
  OAI22XL U4430 ( .A0(n1758), .A1(n3967), .B0(n3186), .B1(n3981), .Y(n2998) );
  OAI22XL U4431 ( .A0(n1759), .A1(n3967), .B0(n3185), .B1(n3981), .Y(n2999) );
  OAI22XL U4432 ( .A0(n1760), .A1(n3967), .B0(n3184), .B1(n3981), .Y(n3000) );
  OAI22XL U4433 ( .A0(n1761), .A1(n3967), .B0(n3183), .B1(n3981), .Y(n3001) );
  OAI22XL U4434 ( .A0(n1762), .A1(n3967), .B0(n3182), .B1(n3981), .Y(n3002) );
  OAI22XL U4435 ( .A0(n1763), .A1(n3967), .B0(n3146), .B1(n3981), .Y(n3003) );
  OAI22XL U4436 ( .A0(n1764), .A1(n3967), .B0(n3145), .B1(n3981), .Y(n3004) );
  OAI22XL U4437 ( .A0(n1765), .A1(n3968), .B0(n3144), .B1(n3981), .Y(n3005) );
  OAI22XL U4438 ( .A0(n1766), .A1(n3968), .B0(n3143), .B1(n3981), .Y(n3006) );
  OAI22XL U4439 ( .A0(n1767), .A1(n3968), .B0(n3142), .B1(n3981), .Y(n3007) );
  OAI22XL U4440 ( .A0(n1768), .A1(n3968), .B0(n3139), .B1(n3982), .Y(n3008) );
  OAI22XL U4441 ( .A0(n1769), .A1(n3968), .B0(n3138), .B1(n3982), .Y(n3009) );
  OAI22XL U4442 ( .A0(n1770), .A1(n3968), .B0(n3137), .B1(n3982), .Y(n3010) );
  OAI22XL U4443 ( .A0(n1771), .A1(n3968), .B0(n3136), .B1(n3982), .Y(n3011) );
  OAI22XL U4444 ( .A0(n1772), .A1(n3968), .B0(n3141), .B1(n3982), .Y(n3012) );
  OAI22XL U4445 ( .A0(n1773), .A1(n3968), .B0(n3135), .B1(n3982), .Y(n3013) );
  OAI22XL U4446 ( .A0(n1774), .A1(n3968), .B0(n3140), .B1(n3982), .Y(n3014) );
  OAI22XL U4447 ( .A0(n1775), .A1(n3968), .B0(n3172), .B1(n3982), .Y(n3015) );
  OAI22XL U4448 ( .A0(n1776), .A1(n3968), .B0(n3180), .B1(n3982), .Y(n3016) );
  OAI22XL U4449 ( .A0(n1777), .A1(n3969), .B0(n3173), .B1(n3982), .Y(n3017) );
  OAI22XL U4450 ( .A0(n1778), .A1(n3969), .B0(n3171), .B1(n3982), .Y(n3018) );
  OAI22XL U4451 ( .A0(n1779), .A1(n3969), .B0(n3189), .B1(n3973), .Y(n3019) );
  OAI22XL U4452 ( .A0(n1780), .A1(n3969), .B0(n3188), .B1(n3984), .Y(n3020) );
  OAI22XL U4453 ( .A0(n1781), .A1(n3969), .B0(n3175), .B1(n3974), .Y(n3021) );
  OAI22XL U4454 ( .A0(n1782), .A1(n3969), .B0(n3181), .B1(n3975), .Y(n3022) );
  OAI22XL U4455 ( .A0(n1783), .A1(n3969), .B0(n3174), .B1(n3978), .Y(n3023) );
  OAI31XL U4456 ( .A0(n3341), .A1(n3313), .A2(n3314), .B0(n430), .Y(n468) );
  AOI22X2 U4457 ( .A0(n3888), .A1(N59), .B0(proc_addr[5]), .B1(n3895), .Y(n181) );
  AOI22X2 U4458 ( .A0(n3888), .A1(N58), .B0(proc_addr[6]), .B1(n3894), .Y(n182) );
  AOI22X2 U4459 ( .A0(n3888), .A1(N57), .B0(proc_addr[7]), .B1(n3897), .Y(n183) );
  AOI22X2 U4460 ( .A0(n3888), .A1(N56), .B0(proc_addr[8]), .B1(n3896), .Y(n184) );
  AOI22X2 U4461 ( .A0(n3888), .A1(N55), .B0(proc_addr[9]), .B1(n3898), .Y(n185) );
  AOI22X2 U4462 ( .A0(n3888), .A1(N54), .B0(proc_addr[10]), .B1(n3899), .Y(
        n186) );
  AOI22X2 U4463 ( .A0(n3888), .A1(N53), .B0(proc_addr[11]), .B1(n3902), .Y(
        n187) );
  AOI22X2 U4464 ( .A0(n3888), .A1(N52), .B0(proc_addr[12]), .B1(n3902), .Y(
        n188) );
  AOI22X2 U4465 ( .A0(n3888), .A1(N51), .B0(proc_addr[13]), .B1(n3902), .Y(
        n189) );
  AOI22X2 U4466 ( .A0(n3888), .A1(N50), .B0(proc_addr[14]), .B1(n3902), .Y(
        n190) );
  AOI22X2 U4467 ( .A0(n3888), .A1(N49), .B0(proc_addr[15]), .B1(n3902), .Y(
        n191) );
  AOI22X2 U4468 ( .A0(n3888), .A1(N48), .B0(proc_addr[16]), .B1(n3902), .Y(
        n192) );
  AOI22X2 U4469 ( .A0(n3888), .A1(N47), .B0(proc_addr[17]), .B1(n3902), .Y(
        n193) );
  AOI22X2 U4470 ( .A0(n3889), .A1(N46), .B0(proc_addr[18]), .B1(n3902), .Y(
        n194) );
  AOI22X2 U4471 ( .A0(n3889), .A1(N45), .B0(proc_addr[19]), .B1(n3900), .Y(
        n195) );
  AOI22X2 U4472 ( .A0(n3889), .A1(N44), .B0(proc_addr[20]), .B1(n3902), .Y(
        n196) );
  AOI22X2 U4473 ( .A0(n3889), .A1(N43), .B0(proc_addr[21]), .B1(n3902), .Y(
        n197) );
  AOI22X2 U4474 ( .A0(n3889), .A1(N42), .B0(proc_addr[22]), .B1(n3902), .Y(
        n198) );
  AOI22X2 U4475 ( .A0(n3889), .A1(N41), .B0(proc_addr[23]), .B1(n3902), .Y(
        n199) );
  AOI22X2 U4476 ( .A0(n3889), .A1(N40), .B0(proc_addr[24]), .B1(n3902), .Y(
        n200) );
  AOI22X2 U4477 ( .A0(n3889), .A1(N38), .B0(proc_addr[26]), .B1(n3901), .Y(
        n202) );
  AOI22X2 U4478 ( .A0(n3889), .A1(N37), .B0(proc_addr[27]), .B1(n3901), .Y(
        n203) );
  AOI22X2 U4479 ( .A0(n3889), .A1(N36), .B0(proc_addr[28]), .B1(n3901), .Y(
        n204) );
  AOI22X2 U4480 ( .A0(n3889), .A1(N35), .B0(proc_addr[29]), .B1(n3901), .Y(
        n205) );
  OAI21XL U4481 ( .A0(n4144), .A1(N34), .B0(n8), .Y(n538) );
  MXI2X1 U4482 ( .A(n3657), .B(n3658), .S0(n3728), .Y(N33) );
  NAND3X2 U4483 ( .A(n3315), .B(n3313), .C(n4143), .Y(n353) );
  OAI22XL U4484 ( .A0(n700), .A1(n3941), .B0(n181), .B1(n3954), .Y(n1940) );
  OAI22XL U4485 ( .A0(n701), .A1(n3941), .B0(n182), .B1(n3954), .Y(n1941) );
  OAI22XL U4486 ( .A0(n702), .A1(n3941), .B0(n183), .B1(n3954), .Y(n1942) );
  OAI22XL U4487 ( .A0(n703), .A1(n3941), .B0(n184), .B1(n3954), .Y(n1943) );
  OAI22XL U4488 ( .A0(n704), .A1(n3942), .B0(n185), .B1(n3954), .Y(n1944) );
  OAI22XL U4489 ( .A0(n705), .A1(n3942), .B0(n186), .B1(n3955), .Y(n1945) );
  OAI22XL U4490 ( .A0(n706), .A1(n3942), .B0(n187), .B1(n3955), .Y(n1946) );
  OAI22XL U4491 ( .A0(n707), .A1(n3942), .B0(n188), .B1(n3955), .Y(n1947) );
  OAI22XL U4492 ( .A0(n708), .A1(n3942), .B0(n189), .B1(n3955), .Y(n1948) );
  OAI22XL U4493 ( .A0(n709), .A1(n3942), .B0(n190), .B1(n3955), .Y(n1949) );
  OAI22XL U4494 ( .A0(n710), .A1(n3942), .B0(n191), .B1(n3955), .Y(n1950) );
  OAI22XL U4495 ( .A0(n711), .A1(n3942), .B0(n192), .B1(n3955), .Y(n1951) );
  OAI22XL U4496 ( .A0(n712), .A1(n3942), .B0(n193), .B1(n3955), .Y(n1952) );
  OAI22XL U4497 ( .A0(n713), .A1(n3942), .B0(n194), .B1(n3955), .Y(n1953) );
  OAI22XL U4498 ( .A0(n714), .A1(n3942), .B0(n195), .B1(n3955), .Y(n1954) );
  OAI22XL U4499 ( .A0(n715), .A1(n3942), .B0(n196), .B1(n3955), .Y(n1955) );
  OAI22XL U4500 ( .A0(n716), .A1(n3943), .B0(n197), .B1(n3956), .Y(n1956) );
  OAI22XL U4501 ( .A0(n717), .A1(n3943), .B0(n198), .B1(n3956), .Y(n1957) );
  OAI22XL U4502 ( .A0(n718), .A1(n3943), .B0(n199), .B1(n3956), .Y(n1958) );
  OAI22XL U4503 ( .A0(n719), .A1(n3943), .B0(n200), .B1(n3956), .Y(n1959) );
  OAI22XL U4504 ( .A0(n720), .A1(n3943), .B0(n201), .B1(n3956), .Y(n1960) );
  OAI22XL U4505 ( .A0(n721), .A1(n3943), .B0(n202), .B1(n3956), .Y(n1961) );
  OAI22XL U4506 ( .A0(n722), .A1(n3943), .B0(n203), .B1(n3956), .Y(n1962) );
  OAI22XL U4507 ( .A0(n723), .A1(n3943), .B0(n204), .B1(n3956), .Y(n1963) );
  OAI22XL U4508 ( .A0(n724), .A1(n3943), .B0(n205), .B1(n3956), .Y(n1964) );
  OAI22XL U4509 ( .A0(n855), .A1(n3913), .B0(n181), .B1(n3923), .Y(n2095) );
  OAI22XL U4510 ( .A0(n856), .A1(n3913), .B0(n182), .B1(n3920), .Y(n2096) );
  OAI22XL U4511 ( .A0(n857), .A1(n3913), .B0(n183), .B1(n3921), .Y(n2097) );
  OAI22XL U4512 ( .A0(n858), .A1(n3913), .B0(n184), .B1(n3916), .Y(n2098) );
  OAI22XL U4513 ( .A0(n859), .A1(n3914), .B0(n185), .B1(n3929), .Y(n2099) );
  OAI22XL U4514 ( .A0(n860), .A1(n3914), .B0(n186), .B1(n3927), .Y(n2100) );
  OAI22XL U4515 ( .A0(n861), .A1(n3914), .B0(n187), .B1(n3927), .Y(n2101) );
  OAI22XL U4516 ( .A0(n862), .A1(n3914), .B0(n188), .B1(n3927), .Y(n2102) );
  OAI22XL U4517 ( .A0(n863), .A1(n3914), .B0(n189), .B1(n3927), .Y(n2103) );
  OAI22XL U4518 ( .A0(n864), .A1(n3914), .B0(n190), .B1(n3927), .Y(n2104) );
  OAI22XL U4519 ( .A0(n865), .A1(n3914), .B0(n191), .B1(n3927), .Y(n2105) );
  OAI22XL U4520 ( .A0(n866), .A1(n3914), .B0(n192), .B1(n3927), .Y(n2106) );
  OAI22XL U4521 ( .A0(n867), .A1(n3914), .B0(n193), .B1(n3927), .Y(n2107) );
  OAI22XL U4522 ( .A0(n868), .A1(n3914), .B0(n194), .B1(n3927), .Y(n2108) );
  OAI22XL U4523 ( .A0(n869), .A1(n3914), .B0(n195), .B1(n3927), .Y(n2109) );
  OAI22XL U4524 ( .A0(n870), .A1(n3914), .B0(n196), .B1(n3927), .Y(n2110) );
  OAI22XL U4525 ( .A0(n871), .A1(n3915), .B0(n197), .B1(n3928), .Y(n2111) );
  OAI22XL U4526 ( .A0(n872), .A1(n3915), .B0(n198), .B1(n3928), .Y(n2112) );
  OAI22XL U4527 ( .A0(n873), .A1(n3915), .B0(n199), .B1(n3928), .Y(n2113) );
  OAI22XL U4528 ( .A0(n874), .A1(n3915), .B0(n200), .B1(n3928), .Y(n2114) );
  OAI22XL U4529 ( .A0(n875), .A1(n3915), .B0(n201), .B1(n3928), .Y(n2115) );
  OAI22XL U4530 ( .A0(n876), .A1(n3915), .B0(n202), .B1(n3928), .Y(n2116) );
  OAI22XL U4531 ( .A0(n877), .A1(n3915), .B0(n203), .B1(n3928), .Y(n2117) );
  OAI22XL U4532 ( .A0(n878), .A1(n3915), .B0(n204), .B1(n3928), .Y(n2118) );
  OAI22XL U4533 ( .A0(n879), .A1(n3915), .B0(n205), .B1(n3928), .Y(n2119) );
  OAI22XL U4534 ( .A0(n1010), .A1(n4099), .B0(n181), .B1(n4113), .Y(n2250) );
  OAI22XL U4535 ( .A0(n1011), .A1(n4099), .B0(n182), .B1(n4111), .Y(n2251) );
  OAI22XL U4536 ( .A0(n1012), .A1(n4099), .B0(n183), .B1(n4112), .Y(n2252) );
  OAI22XL U4537 ( .A0(n1013), .A1(n4099), .B0(n184), .B1(n4112), .Y(n2253) );
  OAI22XL U4538 ( .A0(n1014), .A1(n4099), .B0(n185), .B1(n4112), .Y(n2254) );
  OAI22XL U4539 ( .A0(n1015), .A1(n4099), .B0(n186), .B1(n4112), .Y(n2255) );
  OAI22XL U4540 ( .A0(n1016), .A1(n4099), .B0(n187), .B1(n4112), .Y(n2256) );
  OAI22XL U4541 ( .A0(n1017), .A1(n4099), .B0(n188), .B1(n4112), .Y(n2257) );
  OAI22XL U4542 ( .A0(n1018), .A1(n4099), .B0(n189), .B1(n4112), .Y(n2258) );
  OAI22XL U4543 ( .A0(n1019), .A1(n4099), .B0(n190), .B1(n4112), .Y(n2259) );
  OAI22XL U4544 ( .A0(n1020), .A1(n4100), .B0(n191), .B1(n4113), .Y(n2260) );
  OAI22XL U4545 ( .A0(n1021), .A1(n4100), .B0(n192), .B1(n4113), .Y(n2261) );
  OAI22XL U4546 ( .A0(n1022), .A1(n4100), .B0(n193), .B1(n4113), .Y(n2262) );
  OAI22XL U4547 ( .A0(n1023), .A1(n4100), .B0(n194), .B1(n4113), .Y(n2263) );
  OAI22XL U4548 ( .A0(n1024), .A1(n4100), .B0(n195), .B1(n4113), .Y(n2264) );
  OAI22XL U4549 ( .A0(n1025), .A1(n4100), .B0(n196), .B1(n4113), .Y(n2265) );
  OAI22XL U4550 ( .A0(n1026), .A1(n4100), .B0(n197), .B1(n4113), .Y(n2266) );
  OAI22XL U4551 ( .A0(n1027), .A1(n4100), .B0(n198), .B1(n4113), .Y(n2267) );
  OAI22XL U4552 ( .A0(n1028), .A1(n4100), .B0(n199), .B1(n4113), .Y(n2268) );
  OAI22XL U4553 ( .A0(n1029), .A1(n4100), .B0(n200), .B1(n4113), .Y(n2269) );
  OAI22XL U4554 ( .A0(n1030), .A1(n4100), .B0(n201), .B1(n4113), .Y(n2270) );
  OAI22XL U4555 ( .A0(n1031), .A1(n4100), .B0(n202), .B1(n4114), .Y(n2271) );
  OAI22XL U4556 ( .A0(n1032), .A1(n4101), .B0(n203), .B1(n4114), .Y(n2272) );
  OAI22XL U4557 ( .A0(n1033), .A1(n4101), .B0(n204), .B1(n4114), .Y(n2273) );
  OAI22XL U4558 ( .A0(n1034), .A1(n4101), .B0(n205), .B1(n4114), .Y(n2274) );
  OAI22XL U4559 ( .A0(n1165), .A1(n4081), .B0(n181), .B1(n4091), .Y(n2405) );
  OAI22XL U4560 ( .A0(n1166), .A1(n4081), .B0(n182), .B1(n4088), .Y(n2406) );
  OAI22XL U4561 ( .A0(n1167), .A1(n4081), .B0(n183), .B1(n4089), .Y(n2407) );
  OAI22XL U4562 ( .A0(n1168), .A1(n4081), .B0(n184), .B1(n4084), .Y(n2408) );
  OAI22XL U4563 ( .A0(n1169), .A1(n4082), .B0(n185), .B1(n4097), .Y(n2409) );
  OAI22XL U4564 ( .A0(n1170), .A1(n4082), .B0(n186), .B1(n4095), .Y(n2410) );
  OAI22XL U4565 ( .A0(n1171), .A1(n4082), .B0(n187), .B1(n4095), .Y(n2411) );
  OAI22XL U4566 ( .A0(n1172), .A1(n4082), .B0(n188), .B1(n4095), .Y(n2412) );
  OAI22XL U4567 ( .A0(n1173), .A1(n4082), .B0(n189), .B1(n4095), .Y(n2413) );
  OAI22XL U4568 ( .A0(n1174), .A1(n4082), .B0(n190), .B1(n4095), .Y(n2414) );
  OAI22XL U4569 ( .A0(n1175), .A1(n4082), .B0(n191), .B1(n4095), .Y(n2415) );
  OAI22XL U4570 ( .A0(n1176), .A1(n4082), .B0(n192), .B1(n4095), .Y(n2416) );
  OAI22XL U4571 ( .A0(n1177), .A1(n4082), .B0(n193), .B1(n4095), .Y(n2417) );
  OAI22XL U4572 ( .A0(n1178), .A1(n4082), .B0(n194), .B1(n4095), .Y(n2418) );
  OAI22XL U4573 ( .A0(n1179), .A1(n4082), .B0(n195), .B1(n4095), .Y(n2419) );
  OAI22XL U4574 ( .A0(n1180), .A1(n4082), .B0(n196), .B1(n4095), .Y(n2420) );
  OAI22XL U4575 ( .A0(n1181), .A1(n4083), .B0(n197), .B1(n4096), .Y(n2421) );
  OAI22XL U4576 ( .A0(n1182), .A1(n4083), .B0(n198), .B1(n4096), .Y(n2422) );
  OAI22XL U4577 ( .A0(n1183), .A1(n4083), .B0(n199), .B1(n4096), .Y(n2423) );
  OAI22XL U4578 ( .A0(n1184), .A1(n4083), .B0(n200), .B1(n4096), .Y(n2424) );
  OAI22XL U4579 ( .A0(n1185), .A1(n4083), .B0(n201), .B1(n4096), .Y(n2425) );
  OAI22XL U4580 ( .A0(n1186), .A1(n4083), .B0(n202), .B1(n4096), .Y(n2426) );
  OAI22XL U4581 ( .A0(n1187), .A1(n4083), .B0(n203), .B1(n4096), .Y(n2427) );
  OAI22XL U4582 ( .A0(n1188), .A1(n4083), .B0(n204), .B1(n4096), .Y(n2428) );
  OAI22XL U4583 ( .A0(n1189), .A1(n4083), .B0(n205), .B1(n4096), .Y(n2429) );
  OAI22XL U4584 ( .A0(n1320), .A1(n4053), .B0(n181), .B1(n4066), .Y(n2560) );
  OAI22XL U4585 ( .A0(n1321), .A1(n4053), .B0(n182), .B1(n4066), .Y(n2561) );
  OAI22XL U4586 ( .A0(n1322), .A1(n4053), .B0(n183), .B1(n4066), .Y(n2562) );
  OAI22XL U4587 ( .A0(n1323), .A1(n4053), .B0(n184), .B1(n4066), .Y(n2563) );
  OAI22XL U4588 ( .A0(n1324), .A1(n4054), .B0(n185), .B1(n4066), .Y(n2564) );
  OAI22XL U4589 ( .A0(n1325), .A1(n4054), .B0(n186), .B1(n4067), .Y(n2565) );
  OAI22XL U4590 ( .A0(n1326), .A1(n4054), .B0(n187), .B1(n4067), .Y(n2566) );
  OAI22XL U4591 ( .A0(n1327), .A1(n4054), .B0(n188), .B1(n4067), .Y(n2567) );
  OAI22XL U4592 ( .A0(n1328), .A1(n4054), .B0(n189), .B1(n4067), .Y(n2568) );
  OAI22XL U4593 ( .A0(n1329), .A1(n4054), .B0(n190), .B1(n4067), .Y(n2569) );
  OAI22XL U4594 ( .A0(n1330), .A1(n4054), .B0(n191), .B1(n4067), .Y(n2570) );
  OAI22XL U4595 ( .A0(n1331), .A1(n4054), .B0(n192), .B1(n4067), .Y(n2571) );
  OAI22XL U4596 ( .A0(n1332), .A1(n4054), .B0(n193), .B1(n4067), .Y(n2572) );
  OAI22XL U4597 ( .A0(n1333), .A1(n4054), .B0(n194), .B1(n4067), .Y(n2573) );
  OAI22XL U4598 ( .A0(n1334), .A1(n4054), .B0(n195), .B1(n4067), .Y(n2574) );
  OAI22XL U4599 ( .A0(n1335), .A1(n4054), .B0(n196), .B1(n4067), .Y(n2575) );
  OAI22XL U4600 ( .A0(n1336), .A1(n4048), .B0(n197), .B1(n4068), .Y(n2576) );
  OAI22XL U4601 ( .A0(n1337), .A1(n4046), .B0(n198), .B1(n4068), .Y(n2577) );
  OAI22XL U4602 ( .A0(n1338), .A1(n4044), .B0(n199), .B1(n4068), .Y(n2578) );
  OAI22XL U4603 ( .A0(n1339), .A1(n4043), .B0(n200), .B1(n4068), .Y(n2579) );
  OAI22XL U4604 ( .A0(n1340), .A1(n4048), .B0(n201), .B1(n4068), .Y(n2580) );
  OAI22XL U4605 ( .A0(n1341), .A1(n4046), .B0(n202), .B1(n4068), .Y(n2581) );
  OAI22XL U4606 ( .A0(n1342), .A1(n4044), .B0(n203), .B1(n4068), .Y(n2582) );
  OAI22XL U4607 ( .A0(n1343), .A1(n4043), .B0(n204), .B1(n4068), .Y(n2583) );
  OAI22XL U4608 ( .A0(n1344), .A1(n4043), .B0(n205), .B1(n4068), .Y(n2584) );
  OAI22XL U4609 ( .A0(n1475), .A1(n4025), .B0(n181), .B1(n4035), .Y(n2715) );
  OAI22XL U4610 ( .A0(n1476), .A1(n4025), .B0(n182), .B1(n4032), .Y(n2716) );
  OAI22XL U4611 ( .A0(n1477), .A1(n4025), .B0(n183), .B1(n4033), .Y(n2717) );
  OAI22XL U4612 ( .A0(n1478), .A1(n4025), .B0(n184), .B1(n4028), .Y(n2718) );
  OAI22XL U4613 ( .A0(n1479), .A1(n4026), .B0(n185), .B1(n4041), .Y(n2719) );
  OAI22XL U4614 ( .A0(n1480), .A1(n4026), .B0(n186), .B1(n4039), .Y(n2720) );
  OAI22XL U4615 ( .A0(n1481), .A1(n4026), .B0(n187), .B1(n4039), .Y(n2721) );
  OAI22XL U4616 ( .A0(n1482), .A1(n4026), .B0(n188), .B1(n4039), .Y(n2722) );
  OAI22XL U4617 ( .A0(n1483), .A1(n4026), .B0(n189), .B1(n4039), .Y(n2723) );
  OAI22XL U4618 ( .A0(n1484), .A1(n4026), .B0(n190), .B1(n4039), .Y(n2724) );
  OAI22XL U4619 ( .A0(n1485), .A1(n4026), .B0(n191), .B1(n4039), .Y(n2725) );
  OAI22XL U4620 ( .A0(n1486), .A1(n4026), .B0(n192), .B1(n4039), .Y(n2726) );
  OAI22XL U4621 ( .A0(n1487), .A1(n4026), .B0(n193), .B1(n4039), .Y(n2727) );
  OAI22XL U4622 ( .A0(n1488), .A1(n4026), .B0(n194), .B1(n4039), .Y(n2728) );
  OAI22XL U4623 ( .A0(n1489), .A1(n4026), .B0(n195), .B1(n4039), .Y(n2729) );
  OAI22XL U4624 ( .A0(n1490), .A1(n4026), .B0(n196), .B1(n4039), .Y(n2730) );
  OAI22XL U4625 ( .A0(n1491), .A1(n4027), .B0(n197), .B1(n4040), .Y(n2731) );
  OAI22XL U4626 ( .A0(n1492), .A1(n4027), .B0(n198), .B1(n4040), .Y(n2732) );
  OAI22XL U4627 ( .A0(n1493), .A1(n4027), .B0(n199), .B1(n4040), .Y(n2733) );
  OAI22XL U4628 ( .A0(n1494), .A1(n4027), .B0(n200), .B1(n4040), .Y(n2734) );
  OAI22XL U4629 ( .A0(n1495), .A1(n4027), .B0(n201), .B1(n4040), .Y(n2735) );
  OAI22XL U4630 ( .A0(n1496), .A1(n4027), .B0(n202), .B1(n4040), .Y(n2736) );
  OAI22XL U4631 ( .A0(n1497), .A1(n4027), .B0(n203), .B1(n4040), .Y(n2737) );
  OAI22XL U4632 ( .A0(n1498), .A1(n4027), .B0(n204), .B1(n4040), .Y(n2738) );
  OAI22XL U4633 ( .A0(n1499), .A1(n4027), .B0(n205), .B1(n4040), .Y(n2739) );
  OAI22XL U4634 ( .A0(n1630), .A1(n3997), .B0(n181), .B1(n4010), .Y(n2870) );
  OAI22XL U4635 ( .A0(n1631), .A1(n3997), .B0(n182), .B1(n4010), .Y(n2871) );
  OAI22XL U4636 ( .A0(n1632), .A1(n3997), .B0(n183), .B1(n4010), .Y(n2872) );
  OAI22XL U4637 ( .A0(n1633), .A1(n3997), .B0(n184), .B1(n4010), .Y(n2873) );
  OAI22XL U4638 ( .A0(n1634), .A1(n3998), .B0(n185), .B1(n4010), .Y(n2874) );
  OAI22XL U4639 ( .A0(n1635), .A1(n3998), .B0(n186), .B1(n4011), .Y(n2875) );
  OAI22XL U4640 ( .A0(n1636), .A1(n3998), .B0(n187), .B1(n4011), .Y(n2876) );
  OAI22XL U4641 ( .A0(n1637), .A1(n3998), .B0(n188), .B1(n4011), .Y(n2877) );
  OAI22XL U4642 ( .A0(n1638), .A1(n3998), .B0(n189), .B1(n4011), .Y(n2878) );
  OAI22XL U4643 ( .A0(n1639), .A1(n3998), .B0(n190), .B1(n4011), .Y(n2879) );
  OAI22XL U4644 ( .A0(n1640), .A1(n3998), .B0(n191), .B1(n4011), .Y(n2880) );
  OAI22XL U4645 ( .A0(n1641), .A1(n3998), .B0(n192), .B1(n4011), .Y(n2881) );
  OAI22XL U4646 ( .A0(n1642), .A1(n3998), .B0(n193), .B1(n4011), .Y(n2882) );
  OAI22XL U4647 ( .A0(n1643), .A1(n3998), .B0(n194), .B1(n4011), .Y(n2883) );
  OAI22XL U4648 ( .A0(n1644), .A1(n3998), .B0(n195), .B1(n4011), .Y(n2884) );
  OAI22XL U4649 ( .A0(n1645), .A1(n3998), .B0(n196), .B1(n4011), .Y(n2885) );
  OAI22XL U4650 ( .A0(n1646), .A1(n3992), .B0(n197), .B1(n4012), .Y(n2886) );
  OAI22XL U4651 ( .A0(n1647), .A1(n3990), .B0(n198), .B1(n4012), .Y(n2887) );
  OAI22XL U4652 ( .A0(n1648), .A1(n3988), .B0(n199), .B1(n4012), .Y(n2888) );
  OAI22XL U4653 ( .A0(n1649), .A1(n3987), .B0(n200), .B1(n4012), .Y(n2889) );
  OAI22XL U4654 ( .A0(n1650), .A1(n3992), .B0(n201), .B1(n4012), .Y(n2890) );
  OAI22XL U4655 ( .A0(n1651), .A1(n3990), .B0(n202), .B1(n4012), .Y(n2891) );
  OAI22XL U4656 ( .A0(n1652), .A1(n3988), .B0(n203), .B1(n4012), .Y(n2892) );
  OAI22XL U4657 ( .A0(n1653), .A1(n3987), .B0(n204), .B1(n4012), .Y(n2893) );
  OAI22XL U4658 ( .A0(n1654), .A1(n3987), .B0(n205), .B1(n4012), .Y(n2894) );
  OAI22XL U4659 ( .A0(n1785), .A1(n3969), .B0(n181), .B1(n3979), .Y(n3025) );
  OAI22XL U4660 ( .A0(n1786), .A1(n3969), .B0(n182), .B1(n3976), .Y(n3026) );
  OAI22XL U4661 ( .A0(n1787), .A1(n3969), .B0(n183), .B1(n3977), .Y(n3027) );
  OAI22XL U4662 ( .A0(n1788), .A1(n3969), .B0(n184), .B1(n3972), .Y(n3028) );
  OAI22XL U4663 ( .A0(n1789), .A1(n3970), .B0(n185), .B1(n3985), .Y(n3029) );
  OAI22XL U4664 ( .A0(n1790), .A1(n3970), .B0(n186), .B1(n3983), .Y(n3030) );
  OAI22XL U4665 ( .A0(n1791), .A1(n3970), .B0(n187), .B1(n3983), .Y(n3031) );
  OAI22XL U4666 ( .A0(n1792), .A1(n3970), .B0(n188), .B1(n3983), .Y(n3032) );
  OAI22XL U4667 ( .A0(n1793), .A1(n3970), .B0(n189), .B1(n3983), .Y(n3033) );
  OAI22XL U4668 ( .A0(n1794), .A1(n3970), .B0(n190), .B1(n3983), .Y(n3034) );
  OAI22XL U4669 ( .A0(n1795), .A1(n3970), .B0(n191), .B1(n3983), .Y(n3035) );
  OAI22XL U4670 ( .A0(n1796), .A1(n3970), .B0(n192), .B1(n3983), .Y(n3036) );
  OAI22XL U4671 ( .A0(n1797), .A1(n3970), .B0(n193), .B1(n3983), .Y(n3037) );
  OAI22XL U4672 ( .A0(n1798), .A1(n3970), .B0(n194), .B1(n3983), .Y(n3038) );
  OAI22XL U4673 ( .A0(n1799), .A1(n3970), .B0(n195), .B1(n3983), .Y(n3039) );
  OAI22XL U4674 ( .A0(n1800), .A1(n3970), .B0(n196), .B1(n3983), .Y(n3040) );
  OAI22XL U4675 ( .A0(n1801), .A1(n3971), .B0(n197), .B1(n3984), .Y(n3041) );
  OAI22XL U4676 ( .A0(n1802), .A1(n3971), .B0(n198), .B1(n3984), .Y(n3042) );
  OAI22XL U4677 ( .A0(n1803), .A1(n3971), .B0(n199), .B1(n3984), .Y(n3043) );
  OAI22XL U4678 ( .A0(n1804), .A1(n3971), .B0(n200), .B1(n3984), .Y(n3044) );
  OAI22XL U4679 ( .A0(n1805), .A1(n3971), .B0(n201), .B1(n3984), .Y(n3045) );
  OAI22XL U4680 ( .A0(n1806), .A1(n3971), .B0(n202), .B1(n3984), .Y(n3046) );
  OAI22XL U4681 ( .A0(n1807), .A1(n3971), .B0(n203), .B1(n3984), .Y(n3047) );
  OAI22XL U4682 ( .A0(n1808), .A1(n3971), .B0(n204), .B1(n3984), .Y(n3048) );
  OAI22XL U4683 ( .A0(n1809), .A1(n3971), .B0(n205), .B1(n3984), .Y(n3049) );
  OAI22XL U4684 ( .A0(n725), .A1(n3943), .B0(n206), .B1(n3956), .Y(n1965) );
  OAI22XL U4685 ( .A0(n880), .A1(n3915), .B0(n206), .B1(n3928), .Y(n2120) );
  OAI22XL U4686 ( .A0(n1035), .A1(n4101), .B0(n206), .B1(n4114), .Y(n2275) );
  OAI22XL U4687 ( .A0(n1190), .A1(n4083), .B0(n206), .B1(n4096), .Y(n2430) );
  OAI22XL U4688 ( .A0(n1345), .A1(n4048), .B0(n206), .B1(n4068), .Y(n2585) );
  OAI22XL U4689 ( .A0(n1500), .A1(n4027), .B0(n206), .B1(n4040), .Y(n2740) );
  OAI22XL U4690 ( .A0(n1655), .A1(n3992), .B0(n206), .B1(n4012), .Y(n2895) );
  OAI22XL U4691 ( .A0(n1810), .A1(n3971), .B0(n206), .B1(n3984), .Y(n3050) );
  AND2X2 U4692 ( .A(n534), .B(n3311), .Y(n351) );
  OAI31XL U4693 ( .A0(n7), .A1(N34), .A2(n4144), .B0(n8), .Y(n534) );
  AO22X1 U4694 ( .A0(proc_addr[7]), .A1(mem_read), .B0(N57), .B1(n3872), .Y(
        mem_addr[5]) );
  AO22X1 U4695 ( .A0(proc_addr[10]), .A1(mem_read), .B0(N54), .B1(n3872), .Y(
        mem_addr[8]) );
  AO22X1 U4696 ( .A0(proc_addr[11]), .A1(mem_read), .B0(N53), .B1(n3872), .Y(
        mem_addr[9]) );
  AO22X1 U4697 ( .A0(proc_addr[12]), .A1(mem_read), .B0(N52), .B1(n3872), .Y(
        mem_addr[10]) );
  AO22X1 U4698 ( .A0(proc_addr[17]), .A1(mem_read), .B0(N47), .B1(n3872), .Y(
        mem_addr[15]) );
  AO22X1 U4699 ( .A0(proc_addr[21]), .A1(mem_read), .B0(N43), .B1(n3870), .Y(
        mem_addr[19]) );
  AO22X1 U4700 ( .A0(proc_addr[22]), .A1(mem_read), .B0(N42), .B1(n3872), .Y(
        mem_addr[20]) );
  AO22X1 U4701 ( .A0(proc_addr[23]), .A1(mem_read), .B0(N41), .B1(n3872), .Y(
        mem_addr[21]) );
  AO22X1 U4702 ( .A0(proc_addr[24]), .A1(mem_read), .B0(N40), .B1(mem_write), 
        .Y(mem_addr[22]) );
  AO22X1 U4703 ( .A0(proc_addr[27]), .A1(mem_read), .B0(N37), .B1(n3872), .Y(
        mem_addr[25]) );
  AO22X1 U4704 ( .A0(proc_addr[28]), .A1(mem_read), .B0(N36), .B1(n3872), .Y(
        mem_addr[26]) );
  AO22X1 U4705 ( .A0(proc_addr[29]), .A1(mem_read), .B0(N35), .B1(n3872), .Y(
        mem_addr[27]) );
  AO22X1 U4706 ( .A0(proc_addr[5]), .A1(mem_read), .B0(N59), .B1(n3872), .Y(
        mem_addr[3]) );
  AO22X1 U4707 ( .A0(proc_addr[6]), .A1(mem_read), .B0(N58), .B1(n3872), .Y(
        mem_addr[4]) );
  AO22X1 U4708 ( .A0(proc_addr[8]), .A1(mem_read), .B0(N56), .B1(mem_write), 
        .Y(mem_addr[6]) );
  AO22X1 U4709 ( .A0(proc_addr[9]), .A1(mem_read), .B0(N55), .B1(n3872), .Y(
        mem_addr[7]) );
  AO22X1 U4710 ( .A0(proc_addr[13]), .A1(mem_read), .B0(N51), .B1(n3872), .Y(
        mem_addr[11]) );
  AO22X1 U4711 ( .A0(proc_addr[14]), .A1(mem_read), .B0(N50), .B1(n3872), .Y(
        mem_addr[12]) );
  AO22X1 U4712 ( .A0(proc_addr[15]), .A1(mem_read), .B0(N49), .B1(n3872), .Y(
        mem_addr[13]) );
  AO22X1 U4713 ( .A0(proc_addr[16]), .A1(mem_read), .B0(N48), .B1(n3872), .Y(
        mem_addr[14]) );
  AO22X1 U4714 ( .A0(proc_addr[18]), .A1(mem_read), .B0(N46), .B1(n3872), .Y(
        mem_addr[16]) );
  AO22X1 U4715 ( .A0(proc_addr[19]), .A1(mem_read), .B0(N45), .B1(mem_write), 
        .Y(mem_addr[17]) );
  AO22X1 U4716 ( .A0(proc_addr[20]), .A1(mem_read), .B0(N44), .B1(n3872), .Y(
        mem_addr[18]) );
  AO22X1 U4717 ( .A0(proc_addr[25]), .A1(mem_read), .B0(n3245), .B1(mem_write), 
        .Y(mem_addr[23]) );
  AO22X1 U4718 ( .A0(proc_addr[26]), .A1(mem_read), .B0(N38), .B1(mem_write), 
        .Y(mem_addr[24]) );
  AOI21X2 U4719 ( .A0(n3317), .A1(n3311), .B0(N33), .Y(n207) );
  OAI22XL U4720 ( .A0(n726), .A1(n3943), .B0(n207), .B1(n3956), .Y(n1966) );
  OAI22XL U4721 ( .A0(n881), .A1(n3915), .B0(n207), .B1(n3928), .Y(n2121) );
  OAI22XL U4722 ( .A0(n1036), .A1(n4101), .B0(n207), .B1(n4114), .Y(n2276) );
  OAI22XL U4723 ( .A0(n1191), .A1(n4083), .B0(n207), .B1(n4096), .Y(n2431) );
  OAI22XL U4724 ( .A0(n1346), .A1(n4046), .B0(n207), .B1(n4068), .Y(n2586) );
  OAI22XL U4725 ( .A0(n1501), .A1(n4027), .B0(n207), .B1(n4040), .Y(n2741) );
  OAI22XL U4726 ( .A0(n1656), .A1(n3990), .B0(n207), .B1(n4012), .Y(n2896) );
  OAI22XL U4727 ( .A0(n1811), .A1(n3971), .B0(n207), .B1(n3984), .Y(n3052) );
  MXI4X1 U4728 ( .A(\CACHE[0][64] ), .B(\CACHE[1][64] ), .C(\CACHE[2][64] ), 
        .D(\CACHE[3][64] ), .S0(n3673), .S1(n3704), .Y(n3513) );
  MXI4X1 U4729 ( .A(\CACHE[4][64] ), .B(\CACHE[5][64] ), .C(\CACHE[6][64] ), 
        .D(\CACHE[7][64] ), .S0(n3673), .S1(n3704), .Y(n3514) );
  MXI4X1 U4730 ( .A(\CACHE[0][65] ), .B(\CACHE[1][65] ), .C(\CACHE[2][65] ), 
        .D(\CACHE[3][65] ), .S0(n3673), .S1(n3705), .Y(n3515) );
  MXI4X1 U4731 ( .A(\CACHE[4][65] ), .B(\CACHE[5][65] ), .C(\CACHE[6][65] ), 
        .D(\CACHE[7][65] ), .S0(n3673), .S1(n3705), .Y(n3516) );
  MXI4X1 U4732 ( .A(\CACHE[0][66] ), .B(\CACHE[1][66] ), .C(\CACHE[2][66] ), 
        .D(\CACHE[3][66] ), .S0(n3673), .S1(n3705), .Y(n3517) );
  MXI4X1 U4733 ( .A(\CACHE[4][66] ), .B(\CACHE[5][66] ), .C(\CACHE[6][66] ), 
        .D(\CACHE[7][66] ), .S0(n3673), .S1(n3705), .Y(n3518) );
  MXI4X1 U4734 ( .A(\CACHE[0][67] ), .B(\CACHE[1][67] ), .C(\CACHE[2][67] ), 
        .D(\CACHE[3][67] ), .S0(n3673), .S1(n3705), .Y(n3519) );
  MXI4X1 U4735 ( .A(\CACHE[4][67] ), .B(\CACHE[5][67] ), .C(\CACHE[6][67] ), 
        .D(\CACHE[7][67] ), .S0(n3673), .S1(n3705), .Y(n3520) );
  MXI4X1 U4736 ( .A(\CACHE[0][68] ), .B(\CACHE[1][68] ), .C(\CACHE[2][68] ), 
        .D(\CACHE[3][68] ), .S0(n3673), .S1(n3705), .Y(n3521) );
  MXI4X1 U4737 ( .A(\CACHE[4][68] ), .B(\CACHE[5][68] ), .C(\CACHE[6][68] ), 
        .D(\CACHE[7][68] ), .S0(n3673), .S1(n3705), .Y(n3522) );
  MXI4X1 U4738 ( .A(\CACHE[0][69] ), .B(\CACHE[1][69] ), .C(\CACHE[2][69] ), 
        .D(\CACHE[3][69] ), .S0(n3673), .S1(n3705), .Y(n3523) );
  MXI4X1 U4739 ( .A(\CACHE[4][69] ), .B(\CACHE[5][69] ), .C(\CACHE[6][69] ), 
        .D(\CACHE[7][69] ), .S0(n3673), .S1(n3705), .Y(n3524) );
  MXI4X1 U4740 ( .A(\CACHE[0][70] ), .B(\CACHE[1][70] ), .C(\CACHE[2][70] ), 
        .D(\CACHE[3][70] ), .S0(n3674), .S1(n3705), .Y(n3525) );
  MXI4X1 U4741 ( .A(\CACHE[4][70] ), .B(\CACHE[5][70] ), .C(\CACHE[6][70] ), 
        .D(\CACHE[7][70] ), .S0(n3673), .S1(n3705), .Y(n3526) );
  MXI4X1 U4742 ( .A(\CACHE[0][71] ), .B(\CACHE[1][71] ), .C(\CACHE[2][71] ), 
        .D(\CACHE[3][71] ), .S0(n3674), .S1(n3706), .Y(n3527) );
  MXI4X1 U4743 ( .A(\CACHE[4][71] ), .B(\CACHE[5][71] ), .C(\CACHE[6][71] ), 
        .D(\CACHE[7][71] ), .S0(n3674), .S1(n3706), .Y(n3528) );
  MXI4X1 U4744 ( .A(\CACHE[0][72] ), .B(\CACHE[1][72] ), .C(\CACHE[2][72] ), 
        .D(\CACHE[3][72] ), .S0(n3674), .S1(n3706), .Y(n3529) );
  MXI4X1 U4745 ( .A(\CACHE[4][72] ), .B(\CACHE[5][72] ), .C(\CACHE[6][72] ), 
        .D(\CACHE[7][72] ), .S0(n3674), .S1(n3706), .Y(n3530) );
  MXI4X1 U4746 ( .A(\CACHE[0][73] ), .B(\CACHE[1][73] ), .C(\CACHE[2][73] ), 
        .D(\CACHE[3][73] ), .S0(n3674), .S1(n3706), .Y(n3531) );
  MXI4X1 U4747 ( .A(\CACHE[4][73] ), .B(\CACHE[5][73] ), .C(\CACHE[6][73] ), 
        .D(\CACHE[7][73] ), .S0(n3674), .S1(n3706), .Y(n3532) );
  MXI4X1 U4748 ( .A(\CACHE[0][74] ), .B(\CACHE[1][74] ), .C(\CACHE[2][74] ), 
        .D(\CACHE[3][74] ), .S0(n3674), .S1(n3706), .Y(n3533) );
  MXI4X1 U4749 ( .A(\CACHE[4][74] ), .B(\CACHE[5][74] ), .C(\CACHE[6][74] ), 
        .D(\CACHE[7][74] ), .S0(n3674), .S1(n3706), .Y(n3534) );
  MXI4X1 U4750 ( .A(\CACHE[0][75] ), .B(\CACHE[1][75] ), .C(\CACHE[2][75] ), 
        .D(\CACHE[3][75] ), .S0(n3674), .S1(n3706), .Y(n3535) );
  MXI4X1 U4751 ( .A(\CACHE[4][75] ), .B(\CACHE[5][75] ), .C(\CACHE[6][75] ), 
        .D(\CACHE[7][75] ), .S0(n3674), .S1(n3706), .Y(n3536) );
  MXI4X1 U4752 ( .A(\CACHE[0][76] ), .B(\CACHE[1][76] ), .C(\CACHE[2][76] ), 
        .D(\CACHE[3][76] ), .S0(n3674), .S1(n3706), .Y(n3537) );
  MXI4X1 U4753 ( .A(\CACHE[4][76] ), .B(\CACHE[5][76] ), .C(\CACHE[6][76] ), 
        .D(\CACHE[7][76] ), .S0(n3674), .S1(n3706), .Y(n3538) );
  MXI4X1 U4754 ( .A(\CACHE[0][77] ), .B(\CACHE[1][77] ), .C(\CACHE[2][77] ), 
        .D(\CACHE[3][77] ), .S0(n3675), .S1(n3707), .Y(n3539) );
  MXI4X1 U4755 ( .A(\CACHE[4][77] ), .B(\CACHE[5][77] ), .C(\CACHE[6][77] ), 
        .D(\CACHE[7][77] ), .S0(n3675), .S1(n3707), .Y(n3540) );
  MXI4X1 U4756 ( .A(\CACHE[0][78] ), .B(\CACHE[1][78] ), .C(\CACHE[2][78] ), 
        .D(\CACHE[3][78] ), .S0(n3675), .S1(n3707), .Y(n3541) );
  MXI4X1 U4757 ( .A(\CACHE[4][78] ), .B(\CACHE[5][78] ), .C(\CACHE[6][78] ), 
        .D(\CACHE[7][78] ), .S0(n3675), .S1(n3707), .Y(n3542) );
  MXI4X1 U4758 ( .A(\CACHE[0][79] ), .B(\CACHE[1][79] ), .C(\CACHE[2][79] ), 
        .D(\CACHE[3][79] ), .S0(n3675), .S1(n3707), .Y(n3543) );
  MXI4X1 U4759 ( .A(\CACHE[4][79] ), .B(\CACHE[5][79] ), .C(\CACHE[6][79] ), 
        .D(\CACHE[7][79] ), .S0(n3675), .S1(n3707), .Y(n3544) );
  MXI4X1 U4760 ( .A(\CACHE[0][80] ), .B(\CACHE[1][80] ), .C(\CACHE[2][80] ), 
        .D(\CACHE[3][80] ), .S0(n3675), .S1(n3707), .Y(n3545) );
  MXI4X1 U4761 ( .A(\CACHE[4][80] ), .B(\CACHE[5][80] ), .C(\CACHE[6][80] ), 
        .D(\CACHE[7][80] ), .S0(n3675), .S1(n3707), .Y(n3546) );
  MXI4X1 U4762 ( .A(\CACHE[0][81] ), .B(\CACHE[1][81] ), .C(\CACHE[2][81] ), 
        .D(\CACHE[3][81] ), .S0(n3675), .S1(n3707), .Y(n3547) );
  MXI4X1 U4763 ( .A(\CACHE[4][81] ), .B(\CACHE[5][81] ), .C(\CACHE[6][81] ), 
        .D(\CACHE[7][81] ), .S0(n3675), .S1(n3707), .Y(n3548) );
  MXI4X1 U4764 ( .A(\CACHE[0][82] ), .B(\CACHE[1][82] ), .C(\CACHE[2][82] ), 
        .D(\CACHE[3][82] ), .S0(n3675), .S1(n3707), .Y(n3549) );
  MXI4X1 U4765 ( .A(\CACHE[4][82] ), .B(\CACHE[5][82] ), .C(\CACHE[6][82] ), 
        .D(\CACHE[7][82] ), .S0(n3675), .S1(n3707), .Y(n3550) );
  MXI4X1 U4766 ( .A(\CACHE[0][83] ), .B(\CACHE[1][83] ), .C(\CACHE[2][83] ), 
        .D(\CACHE[3][83] ), .S0(n3676), .S1(n3709), .Y(n3551) );
  MXI4X1 U4767 ( .A(\CACHE[4][83] ), .B(\CACHE[5][83] ), .C(\CACHE[6][83] ), 
        .D(\CACHE[7][83] ), .S0(n3675), .S1(n3710), .Y(n3552) );
  MXI4X1 U4768 ( .A(\CACHE[0][84] ), .B(\CACHE[1][84] ), .C(\CACHE[2][84] ), 
        .D(\CACHE[3][84] ), .S0(n3676), .S1(n3693), .Y(n3553) );
  MXI4X1 U4769 ( .A(\CACHE[4][84] ), .B(\CACHE[5][84] ), .C(\CACHE[6][84] ), 
        .D(\CACHE[7][84] ), .S0(n3676), .S1(n3694), .Y(n3554) );
  MXI4X1 U4770 ( .A(\CACHE[0][85] ), .B(\CACHE[1][85] ), .C(\CACHE[2][85] ), 
        .D(\CACHE[3][85] ), .S0(n3676), .S1(n3687), .Y(n3555) );
  MXI4X1 U4771 ( .A(\CACHE[4][85] ), .B(\CACHE[5][85] ), .C(\CACHE[6][85] ), 
        .D(\CACHE[7][85] ), .S0(n3676), .S1(n3694), .Y(n3556) );
  MXI4X1 U4772 ( .A(\CACHE[0][86] ), .B(\CACHE[1][86] ), .C(\CACHE[2][86] ), 
        .D(\CACHE[3][86] ), .S0(n3676), .S1(n3700), .Y(n3557) );
  MXI4X1 U4773 ( .A(\CACHE[4][86] ), .B(\CACHE[5][86] ), .C(\CACHE[6][86] ), 
        .D(\CACHE[7][86] ), .S0(n3676), .S1(n3697), .Y(n3558) );
  MXI4X1 U4774 ( .A(\CACHE[0][87] ), .B(\CACHE[1][87] ), .C(\CACHE[2][87] ), 
        .D(\CACHE[3][87] ), .S0(n3676), .S1(n3686), .Y(n3559) );
  MXI4X1 U4775 ( .A(\CACHE[4][87] ), .B(\CACHE[5][87] ), .C(\CACHE[6][87] ), 
        .D(\CACHE[7][87] ), .S0(n3676), .S1(n3708), .Y(n3560) );
  MXI4X1 U4776 ( .A(\CACHE[0][88] ), .B(\CACHE[1][88] ), .C(\CACHE[2][88] ), 
        .D(\CACHE[3][88] ), .S0(n3676), .S1(n3697), .Y(n3561) );
  MXI4X1 U4777 ( .A(\CACHE[4][88] ), .B(\CACHE[5][88] ), .C(\CACHE[6][88] ), 
        .D(\CACHE[7][88] ), .S0(n3676), .S1(n3699), .Y(n3562) );
  MXI4X1 U4778 ( .A(\CACHE[0][89] ), .B(\CACHE[1][89] ), .C(\CACHE[2][89] ), 
        .D(\CACHE[3][89] ), .S0(n3676), .S1(n3707), .Y(n3563) );
  MXI4X1 U4779 ( .A(\CACHE[4][89] ), .B(\CACHE[5][89] ), .C(\CACHE[6][89] ), 
        .D(\CACHE[7][89] ), .S0(n3676), .S1(n3707), .Y(n3564) );
  MXI4X1 U4780 ( .A(\CACHE[0][90] ), .B(\CACHE[1][90] ), .C(\CACHE[2][90] ), 
        .D(\CACHE[3][90] ), .S0(n3677), .S1(n3698), .Y(n3565) );
  MXI4X1 U4781 ( .A(\CACHE[4][90] ), .B(\CACHE[5][90] ), .C(\CACHE[6][90] ), 
        .D(\CACHE[7][90] ), .S0(n3677), .S1(n3698), .Y(n3566) );
  MXI4X1 U4782 ( .A(\CACHE[0][91] ), .B(\CACHE[1][91] ), .C(\CACHE[2][91] ), 
        .D(\CACHE[3][91] ), .S0(n3677), .S1(n3701), .Y(n3567) );
  MXI4X1 U4783 ( .A(\CACHE[4][91] ), .B(\CACHE[5][91] ), .C(\CACHE[6][91] ), 
        .D(\CACHE[7][91] ), .S0(n3677), .S1(n3701), .Y(n3568) );
  MXI4X1 U4784 ( .A(\CACHE[0][92] ), .B(\CACHE[1][92] ), .C(\CACHE[2][92] ), 
        .D(\CACHE[3][92] ), .S0(n3677), .S1(n3703), .Y(n3569) );
  MXI4X1 U4785 ( .A(\CACHE[4][92] ), .B(\CACHE[5][92] ), .C(\CACHE[6][92] ), 
        .D(\CACHE[7][92] ), .S0(n3677), .S1(n3703), .Y(n3570) );
  MXI4X1 U4786 ( .A(\CACHE[0][93] ), .B(\CACHE[1][93] ), .C(\CACHE[2][93] ), 
        .D(\CACHE[3][93] ), .S0(n3677), .S1(n3704), .Y(n3571) );
  MXI4X1 U4787 ( .A(\CACHE[4][93] ), .B(\CACHE[5][93] ), .C(\CACHE[6][93] ), 
        .D(\CACHE[7][93] ), .S0(n3677), .S1(n3701), .Y(n3572) );
  MXI4X1 U4788 ( .A(\CACHE[0][94] ), .B(\CACHE[1][94] ), .C(\CACHE[2][94] ), 
        .D(\CACHE[3][94] ), .S0(n3677), .S1(n3705), .Y(n3573) );
  MXI4X1 U4789 ( .A(\CACHE[4][94] ), .B(\CACHE[5][94] ), .C(\CACHE[6][94] ), 
        .D(\CACHE[7][94] ), .S0(n3677), .S1(n3703), .Y(n3574) );
  MXI4X1 U4790 ( .A(\CACHE[0][95] ), .B(\CACHE[1][95] ), .C(\CACHE[2][95] ), 
        .D(\CACHE[3][95] ), .S0(n3677), .S1(n3708), .Y(n3575) );
  MXI4X1 U4791 ( .A(\CACHE[4][95] ), .B(\CACHE[5][95] ), .C(\CACHE[6][95] ), 
        .D(\CACHE[7][95] ), .S0(n3677), .S1(n3708), .Y(n3576) );
  MXI4X1 U4792 ( .A(\CACHE[0][32] ), .B(\CACHE[1][32] ), .C(\CACHE[2][32] ), 
        .D(\CACHE[3][32] ), .S0(n3669), .S1(n3700), .Y(n3449) );
  MXI4X1 U4793 ( .A(\CACHE[4][32] ), .B(\CACHE[5][32] ), .C(\CACHE[6][32] ), 
        .D(\CACHE[7][32] ), .S0(n3669), .S1(n3700), .Y(n3450) );
  MXI4X1 U4794 ( .A(\CACHE[0][33] ), .B(\CACHE[1][33] ), .C(\CACHE[2][33] ), 
        .D(\CACHE[3][33] ), .S0(n3669), .S1(n3700), .Y(n3451) );
  MXI4X1 U4795 ( .A(\CACHE[4][33] ), .B(\CACHE[5][33] ), .C(\CACHE[6][33] ), 
        .D(\CACHE[7][33] ), .S0(n3669), .S1(n3700), .Y(n3452) );
  MXI4X1 U4796 ( .A(\CACHE[0][34] ), .B(\CACHE[1][34] ), .C(\CACHE[2][34] ), 
        .D(\CACHE[3][34] ), .S0(n3669), .S1(n3700), .Y(n3453) );
  MXI4X1 U4797 ( .A(\CACHE[4][34] ), .B(\CACHE[5][34] ), .C(\CACHE[6][34] ), 
        .D(\CACHE[7][34] ), .S0(n3669), .S1(n3700), .Y(n3454) );
  MXI4X1 U4798 ( .A(\CACHE[0][35] ), .B(\CACHE[1][35] ), .C(\CACHE[2][35] ), 
        .D(\CACHE[3][35] ), .S0(n3669), .S1(n3701), .Y(n3455) );
  MXI4X1 U4799 ( .A(\CACHE[4][35] ), .B(\CACHE[5][35] ), .C(\CACHE[6][35] ), 
        .D(\CACHE[7][35] ), .S0(n3669), .S1(n3701), .Y(n3456) );
  MXI4X1 U4800 ( .A(\CACHE[0][36] ), .B(\CACHE[1][36] ), .C(\CACHE[2][36] ), 
        .D(\CACHE[3][36] ), .S0(n3669), .S1(n3701), .Y(n3457) );
  MXI4X1 U4801 ( .A(\CACHE[4][36] ), .B(\CACHE[5][36] ), .C(\CACHE[6][36] ), 
        .D(\CACHE[7][36] ), .S0(n3669), .S1(n3701), .Y(n3458) );
  MXI4X1 U4802 ( .A(\CACHE[0][37] ), .B(\CACHE[1][37] ), .C(\CACHE[2][37] ), 
        .D(\CACHE[3][37] ), .S0(n3669), .S1(n3701), .Y(n3459) );
  MXI4X1 U4803 ( .A(\CACHE[4][37] ), .B(\CACHE[5][37] ), .C(\CACHE[6][37] ), 
        .D(\CACHE[7][37] ), .S0(n3669), .S1(n3701), .Y(n3460) );
  MXI4X1 U4804 ( .A(\CACHE[0][38] ), .B(\CACHE[1][38] ), .C(\CACHE[2][38] ), 
        .D(\CACHE[3][38] ), .S0(n3670), .S1(n3701), .Y(n3461) );
  MXI4X1 U4805 ( .A(\CACHE[4][38] ), .B(\CACHE[5][38] ), .C(\CACHE[6][38] ), 
        .D(\CACHE[7][38] ), .S0(n3670), .S1(n3701), .Y(n3462) );
  MXI4X1 U4806 ( .A(\CACHE[0][39] ), .B(\CACHE[1][39] ), .C(\CACHE[2][39] ), 
        .D(\CACHE[3][39] ), .S0(n3670), .S1(n3701), .Y(n3463) );
  MXI4X1 U4807 ( .A(\CACHE[4][39] ), .B(\CACHE[5][39] ), .C(\CACHE[6][39] ), 
        .D(\CACHE[7][39] ), .S0(n3670), .S1(n3701), .Y(n3464) );
  MXI4X1 U4808 ( .A(\CACHE[0][40] ), .B(\CACHE[1][40] ), .C(\CACHE[2][40] ), 
        .D(\CACHE[3][40] ), .S0(n3670), .S1(n3701), .Y(n3465) );
  MXI4X1 U4809 ( .A(\CACHE[4][40] ), .B(\CACHE[5][40] ), .C(\CACHE[6][40] ), 
        .D(\CACHE[7][40] ), .S0(n3670), .S1(n3701), .Y(n3466) );
  MXI4X1 U4810 ( .A(\CACHE[0][41] ), .B(\CACHE[1][41] ), .C(\CACHE[2][41] ), 
        .D(\CACHE[3][41] ), .S0(n3670), .S1(n3702), .Y(n3467) );
  MXI4X1 U4811 ( .A(\CACHE[4][41] ), .B(\CACHE[5][41] ), .C(\CACHE[6][41] ), 
        .D(\CACHE[7][41] ), .S0(n3670), .S1(n3702), .Y(n3468) );
  MXI4X1 U4812 ( .A(\CACHE[0][42] ), .B(\CACHE[1][42] ), .C(\CACHE[2][42] ), 
        .D(\CACHE[3][42] ), .S0(n3670), .S1(n3702), .Y(n3469) );
  MXI4X1 U4813 ( .A(\CACHE[4][42] ), .B(\CACHE[5][42] ), .C(\CACHE[6][42] ), 
        .D(\CACHE[7][42] ), .S0(n3670), .S1(n3702), .Y(n3470) );
  MXI4X1 U4814 ( .A(\CACHE[0][43] ), .B(\CACHE[1][43] ), .C(\CACHE[2][43] ), 
        .D(\CACHE[3][43] ), .S0(n3670), .S1(n3702), .Y(n3471) );
  MXI4X1 U4815 ( .A(\CACHE[4][43] ), .B(\CACHE[5][43] ), .C(\CACHE[6][43] ), 
        .D(\CACHE[7][43] ), .S0(n3670), .S1(n3702), .Y(n3472) );
  MXI4X1 U4816 ( .A(\CACHE[0][44] ), .B(\CACHE[1][44] ), .C(\CACHE[2][44] ), 
        .D(\CACHE[3][44] ), .S0(n3671), .S1(n3702), .Y(n3473) );
  MXI4X1 U4817 ( .A(\CACHE[4][44] ), .B(\CACHE[5][44] ), .C(\CACHE[6][44] ), 
        .D(\CACHE[7][44] ), .S0(n3670), .S1(n3702), .Y(n3474) );
  MXI4X1 U4818 ( .A(\CACHE[0][45] ), .B(\CACHE[1][45] ), .C(\CACHE[2][45] ), 
        .D(\CACHE[3][45] ), .S0(n3671), .S1(n3702), .Y(n3475) );
  MXI4X1 U4819 ( .A(\CACHE[4][45] ), .B(\CACHE[5][45] ), .C(\CACHE[6][45] ), 
        .D(\CACHE[7][45] ), .S0(n3671), .S1(n3702), .Y(n3476) );
  MXI4X1 U4820 ( .A(\CACHE[0][46] ), .B(\CACHE[1][46] ), .C(\CACHE[2][46] ), 
        .D(\CACHE[3][46] ), .S0(n3671), .S1(n3702), .Y(n3477) );
  MXI4X1 U4821 ( .A(\CACHE[4][46] ), .B(\CACHE[5][46] ), .C(\CACHE[6][46] ), 
        .D(\CACHE[7][46] ), .S0(n3671), .S1(n3702), .Y(n3478) );
  MXI4X1 U4822 ( .A(\CACHE[0][47] ), .B(\CACHE[1][47] ), .C(\CACHE[2][47] ), 
        .D(\CACHE[3][47] ), .S0(n3671), .S1(n3703), .Y(n3479) );
  MXI4X1 U4823 ( .A(\CACHE[4][47] ), .B(\CACHE[5][47] ), .C(\CACHE[6][47] ), 
        .D(\CACHE[7][47] ), .S0(n3671), .S1(n3703), .Y(n3480) );
  MXI4X1 U4824 ( .A(\CACHE[0][48] ), .B(\CACHE[1][48] ), .C(\CACHE[2][48] ), 
        .D(\CACHE[3][48] ), .S0(n3671), .S1(n3703), .Y(n3481) );
  MXI4X1 U4825 ( .A(\CACHE[4][48] ), .B(\CACHE[5][48] ), .C(\CACHE[6][48] ), 
        .D(\CACHE[7][48] ), .S0(n3671), .S1(n3703), .Y(n3482) );
  MXI4X1 U4826 ( .A(\CACHE[0][49] ), .B(\CACHE[1][49] ), .C(\CACHE[2][49] ), 
        .D(\CACHE[3][49] ), .S0(n3671), .S1(n3703), .Y(n3483) );
  MXI4X1 U4827 ( .A(\CACHE[4][49] ), .B(\CACHE[5][49] ), .C(\CACHE[6][49] ), 
        .D(\CACHE[7][49] ), .S0(n3671), .S1(n3703), .Y(n3484) );
  MXI4X1 U4828 ( .A(\CACHE[0][50] ), .B(\CACHE[1][50] ), .C(\CACHE[2][50] ), 
        .D(\CACHE[3][50] ), .S0(n3671), .S1(n3703), .Y(n3485) );
  MXI4X1 U4829 ( .A(\CACHE[4][50] ), .B(\CACHE[5][50] ), .C(\CACHE[6][50] ), 
        .D(\CACHE[7][50] ), .S0(n3671), .S1(n3703), .Y(n3486) );
  MXI4X1 U4830 ( .A(\CACHE[0][51] ), .B(\CACHE[1][51] ), .C(\CACHE[2][51] ), 
        .D(\CACHE[3][51] ), .S0(n3665), .S1(n3703), .Y(n3487) );
  MXI4X1 U4831 ( .A(\CACHE[4][51] ), .B(\CACHE[5][51] ), .C(\CACHE[6][51] ), 
        .D(\CACHE[7][51] ), .S0(n3679), .S1(n3703), .Y(n3488) );
  MXI4X1 U4832 ( .A(\CACHE[0][52] ), .B(\CACHE[1][52] ), .C(\CACHE[2][52] ), 
        .D(\CACHE[3][52] ), .S0(n3664), .S1(n3703), .Y(n3489) );
  MXI4X1 U4833 ( .A(\CACHE[4][52] ), .B(\CACHE[5][52] ), .C(\CACHE[6][52] ), 
        .D(\CACHE[7][52] ), .S0(n3674), .S1(n3703), .Y(n3490) );
  MXI4X1 U4834 ( .A(\CACHE[0][53] ), .B(\CACHE[1][53] ), .C(\CACHE[2][53] ), 
        .D(\CACHE[3][53] ), .S0(n3669), .S1(n3700), .Y(n3491) );
  MXI4X1 U4835 ( .A(\CACHE[4][53] ), .B(\CACHE[5][53] ), .C(\CACHE[6][53] ), 
        .D(\CACHE[7][53] ), .S0(n3680), .S1(n3699), .Y(n3492) );
  MXI4X1 U4836 ( .A(\CACHE[0][54] ), .B(\CACHE[1][54] ), .C(\CACHE[2][54] ), 
        .D(\CACHE[3][54] ), .S0(n3673), .S1(n3696), .Y(n3493) );
  MXI4X1 U4837 ( .A(\CACHE[4][54] ), .B(\CACHE[5][54] ), .C(\CACHE[6][54] ), 
        .D(\CACHE[7][54] ), .S0(n3666), .S1(n3710), .Y(n3494) );
  MXI4X1 U4838 ( .A(\CACHE[0][55] ), .B(\CACHE[1][55] ), .C(\CACHE[2][55] ), 
        .D(\CACHE[3][55] ), .S0(n3671), .S1(n3699), .Y(n3495) );
  MXI4X1 U4839 ( .A(\CACHE[4][55] ), .B(\CACHE[5][55] ), .C(\CACHE[6][55] ), 
        .D(\CACHE[7][55] ), .S0(n3676), .S1(n3703), .Y(n3496) );
  MXI4X1 U4840 ( .A(\CACHE[0][56] ), .B(\CACHE[1][56] ), .C(\CACHE[2][56] ), 
        .D(\CACHE[3][56] ), .S0(n3668), .S1(n3710), .Y(n3497) );
  MXI4X1 U4841 ( .A(\CACHE[4][56] ), .B(\CACHE[5][56] ), .C(\CACHE[6][56] ), 
        .D(\CACHE[7][56] ), .S0(n3675), .S1(n3701), .Y(n3498) );
  MXI4X1 U4842 ( .A(\CACHE[0][57] ), .B(\CACHE[1][57] ), .C(\CACHE[2][57] ), 
        .D(\CACHE[3][57] ), .S0(n3672), .S1(n3700), .Y(n3499) );
  MXI4X1 U4843 ( .A(\CACHE[4][57] ), .B(\CACHE[5][57] ), .C(\CACHE[6][57] ), 
        .D(\CACHE[7][57] ), .S0(n3670), .S1(n3702), .Y(n3500) );
  MXI4X1 U4844 ( .A(\CACHE[0][58] ), .B(\CACHE[1][58] ), .C(\CACHE[2][58] ), 
        .D(\CACHE[3][58] ), .S0(n3672), .S1(n3704), .Y(n3501) );
  MXI4X1 U4845 ( .A(\CACHE[4][58] ), .B(\CACHE[5][58] ), .C(\CACHE[6][58] ), 
        .D(\CACHE[7][58] ), .S0(n3672), .S1(n3705), .Y(n3502) );
  MXI4X1 U4846 ( .A(\CACHE[0][59] ), .B(\CACHE[1][59] ), .C(\CACHE[2][59] ), 
        .D(\CACHE[3][59] ), .S0(n3672), .S1(n3704), .Y(n3503) );
  MXI4X1 U4847 ( .A(\CACHE[4][59] ), .B(\CACHE[5][59] ), .C(\CACHE[6][59] ), 
        .D(\CACHE[7][59] ), .S0(n3672), .S1(n3704), .Y(n3504) );
  MXI4X1 U4848 ( .A(\CACHE[0][60] ), .B(\CACHE[1][60] ), .C(\CACHE[2][60] ), 
        .D(\CACHE[3][60] ), .S0(n3672), .S1(n3704), .Y(n3505) );
  MXI4X1 U4849 ( .A(\CACHE[4][60] ), .B(\CACHE[5][60] ), .C(\CACHE[6][60] ), 
        .D(\CACHE[7][60] ), .S0(n3672), .S1(n3704), .Y(n3506) );
  MXI4X1 U4850 ( .A(\CACHE[0][61] ), .B(\CACHE[1][61] ), .C(\CACHE[2][61] ), 
        .D(\CACHE[3][61] ), .S0(n3672), .S1(n3704), .Y(n3507) );
  MXI4X1 U4851 ( .A(\CACHE[4][61] ), .B(\CACHE[5][61] ), .C(\CACHE[6][61] ), 
        .D(\CACHE[7][61] ), .S0(n3672), .S1(n3704), .Y(n3508) );
  MXI4X1 U4852 ( .A(\CACHE[0][62] ), .B(\CACHE[1][62] ), .C(\CACHE[2][62] ), 
        .D(\CACHE[3][62] ), .S0(n3672), .S1(n3704), .Y(n3509) );
  MXI4X1 U4853 ( .A(\CACHE[4][62] ), .B(\CACHE[5][62] ), .C(\CACHE[6][62] ), 
        .D(\CACHE[7][62] ), .S0(n3672), .S1(n3704), .Y(n3510) );
  MXI4X1 U4854 ( .A(\CACHE[0][63] ), .B(\CACHE[1][63] ), .C(\CACHE[2][63] ), 
        .D(\CACHE[3][63] ), .S0(n3672), .S1(n3704), .Y(n3511) );
  MXI4X1 U4855 ( .A(\CACHE[4][63] ), .B(\CACHE[5][63] ), .C(\CACHE[6][63] ), 
        .D(\CACHE[7][63] ), .S0(n3672), .S1(n3704), .Y(n3512) );
  MXI4X1 U4856 ( .A(\CACHE[0][0] ), .B(\CACHE[1][0] ), .C(\CACHE[2][0] ), .D(
        \CACHE[3][0] ), .S0(n3665), .S1(n3696), .Y(n3385) );
  MXI4X1 U4857 ( .A(\CACHE[4][0] ), .B(\CACHE[5][0] ), .C(\CACHE[6][0] ), .D(
        \CACHE[7][0] ), .S0(n3665), .S1(n3696), .Y(n3386) );
  MXI4X1 U4858 ( .A(\CACHE[0][1] ), .B(\CACHE[1][1] ), .C(\CACHE[2][1] ), .D(
        \CACHE[3][1] ), .S0(n3665), .S1(n3696), .Y(n3387) );
  MXI4X1 U4859 ( .A(\CACHE[4][1] ), .B(\CACHE[5][1] ), .C(\CACHE[6][1] ), .D(
        \CACHE[7][1] ), .S0(n3665), .S1(n3696), .Y(n3388) );
  MXI4X1 U4860 ( .A(\CACHE[0][2] ), .B(\CACHE[1][2] ), .C(\CACHE[2][2] ), .D(
        \CACHE[3][2] ), .S0(n3665), .S1(n3696), .Y(n3389) );
  MXI4X1 U4861 ( .A(\CACHE[4][2] ), .B(\CACHE[5][2] ), .C(\CACHE[6][2] ), .D(
        \CACHE[7][2] ), .S0(n3665), .S1(n3696), .Y(n3390) );
  MXI4X1 U4862 ( .A(\CACHE[0][3] ), .B(\CACHE[1][3] ), .C(\CACHE[2][3] ), .D(
        \CACHE[3][3] ), .S0(n3665), .S1(n3696), .Y(n3391) );
  MXI4X1 U4863 ( .A(\CACHE[4][3] ), .B(\CACHE[5][3] ), .C(\CACHE[6][3] ), .D(
        \CACHE[7][3] ), .S0(n3665), .S1(n3696), .Y(n3392) );
  MXI4X1 U4864 ( .A(\CACHE[0][4] ), .B(\CACHE[1][4] ), .C(\CACHE[2][4] ), .D(
        \CACHE[3][4] ), .S0(n3665), .S1(n3696), .Y(n3393) );
  MXI4X1 U4865 ( .A(\CACHE[4][4] ), .B(\CACHE[5][4] ), .C(\CACHE[6][4] ), .D(
        \CACHE[7][4] ), .S0(n3665), .S1(n3696), .Y(n3394) );
  MXI4X1 U4866 ( .A(\CACHE[4][5] ), .B(\CACHE[5][5] ), .C(\CACHE[6][5] ), .D(
        \CACHE[7][5] ), .S0(n3665), .S1(n3697), .Y(n3396) );
  MXI4X1 U4867 ( .A(\CACHE[0][5] ), .B(\CACHE[1][5] ), .C(\CACHE[2][5] ), .D(
        \CACHE[3][5] ), .S0(n3677), .S1(n3697), .Y(n3395) );
  MXI4X1 U4868 ( .A(\CACHE[0][6] ), .B(\CACHE[1][6] ), .C(\CACHE[2][6] ), .D(
        \CACHE[3][6] ), .S0(n3672), .S1(n3697), .Y(n3397) );
  MXI4X1 U4869 ( .A(\CACHE[4][6] ), .B(\CACHE[5][6] ), .C(\CACHE[6][6] ), .D(
        \CACHE[7][6] ), .S0(n3674), .S1(n3697), .Y(n3398) );
  MXI4X1 U4870 ( .A(\CACHE[0][7] ), .B(\CACHE[1][7] ), .C(\CACHE[2][7] ), .D(
        \CACHE[3][7] ), .S0(n3678), .S1(n3697), .Y(n3399) );
  MXI4X1 U4871 ( .A(\CACHE[4][7] ), .B(\CACHE[5][7] ), .C(\CACHE[6][7] ), .D(
        \CACHE[7][7] ), .S0(n3667), .S1(n3697), .Y(n3400) );
  MXI4X1 U4872 ( .A(\CACHE[0][8] ), .B(\CACHE[1][8] ), .C(\CACHE[2][8] ), .D(
        \CACHE[3][8] ), .S0(n3675), .S1(n3697), .Y(n3401) );
  MXI4X1 U4873 ( .A(\CACHE[4][8] ), .B(\CACHE[5][8] ), .C(\CACHE[6][8] ), .D(
        \CACHE[7][8] ), .S0(n3678), .S1(n3697), .Y(n3402) );
  MXI4X1 U4874 ( .A(\CACHE[0][9] ), .B(\CACHE[1][9] ), .C(\CACHE[2][9] ), .D(
        \CACHE[3][9] ), .S0(n3670), .S1(n3697), .Y(n3403) );
  MXI4X1 U4875 ( .A(\CACHE[4][9] ), .B(\CACHE[5][9] ), .C(\CACHE[6][9] ), .D(
        \CACHE[7][9] ), .S0(n3677), .S1(n3697), .Y(n3404) );
  MXI4X1 U4876 ( .A(\CACHE[0][10] ), .B(\CACHE[1][10] ), .C(\CACHE[2][10] ), 
        .D(\CACHE[3][10] ), .S0(n3669), .S1(n3697), .Y(n3405) );
  MXI4X1 U4877 ( .A(\CACHE[4][10] ), .B(\CACHE[5][10] ), .C(\CACHE[6][10] ), 
        .D(\CACHE[7][10] ), .S0(n3672), .S1(n3697), .Y(n3406) );
  MXI4X1 U4878 ( .A(\CACHE[0][11] ), .B(\CACHE[1][11] ), .C(\CACHE[2][11] ), 
        .D(\CACHE[3][11] ), .S0(n3667), .S1(n3698), .Y(n3407) );
  MXI4X1 U4879 ( .A(\CACHE[4][11] ), .B(\CACHE[5][11] ), .C(\CACHE[6][11] ), 
        .D(\CACHE[7][11] ), .S0(n3676), .S1(n3698), .Y(n3408) );
  MXI4X1 U4880 ( .A(\CACHE[0][12] ), .B(\CACHE[1][12] ), .C(\CACHE[2][12] ), 
        .D(\CACHE[3][12] ), .S0(n3666), .S1(n3698), .Y(n3409) );
  MXI4X1 U4881 ( .A(\CACHE[4][12] ), .B(\CACHE[5][12] ), .C(\CACHE[6][12] ), 
        .D(\CACHE[7][12] ), .S0(n3666), .S1(n3698), .Y(n3410) );
  MXI4X1 U4882 ( .A(\CACHE[0][13] ), .B(\CACHE[1][13] ), .C(\CACHE[2][13] ), 
        .D(\CACHE[3][13] ), .S0(n3666), .S1(n3698), .Y(n3411) );
  MXI4X1 U4883 ( .A(\CACHE[4][13] ), .B(\CACHE[5][13] ), .C(\CACHE[6][13] ), 
        .D(\CACHE[7][13] ), .S0(n3666), .S1(n3698), .Y(n3412) );
  MXI4X1 U4884 ( .A(\CACHE[0][14] ), .B(\CACHE[1][14] ), .C(\CACHE[2][14] ), 
        .D(\CACHE[3][14] ), .S0(n3666), .S1(n3698), .Y(n3413) );
  MXI4X1 U4885 ( .A(\CACHE[4][14] ), .B(\CACHE[5][14] ), .C(\CACHE[6][14] ), 
        .D(\CACHE[7][14] ), .S0(n3666), .S1(n3698), .Y(n3414) );
  MXI4X1 U4886 ( .A(\CACHE[0][15] ), .B(\CACHE[1][15] ), .C(\CACHE[2][15] ), 
        .D(\CACHE[3][15] ), .S0(n3666), .S1(n3698), .Y(n3415) );
  MXI4X1 U4887 ( .A(\CACHE[4][15] ), .B(\CACHE[5][15] ), .C(\CACHE[6][15] ), 
        .D(\CACHE[7][15] ), .S0(n3666), .S1(n3698), .Y(n3416) );
  MXI4X1 U4888 ( .A(\CACHE[0][16] ), .B(\CACHE[1][16] ), .C(\CACHE[2][16] ), 
        .D(\CACHE[3][16] ), .S0(n3666), .S1(n3698), .Y(n3417) );
  MXI4X1 U4889 ( .A(\CACHE[4][16] ), .B(\CACHE[5][16] ), .C(\CACHE[6][16] ), 
        .D(\CACHE[7][16] ), .S0(n3666), .S1(n3698), .Y(n3418) );
  MXI4X1 U4890 ( .A(\CACHE[0][17] ), .B(\CACHE[1][17] ), .C(\CACHE[2][17] ), 
        .D(\CACHE[3][17] ), .S0(n3666), .S1(n3697), .Y(n3419) );
  MXI4X1 U4891 ( .A(\CACHE[4][17] ), .B(\CACHE[5][17] ), .C(\CACHE[6][17] ), 
        .D(\CACHE[7][17] ), .S0(n3666), .S1(n3686), .Y(n3420) );
  MXI4X1 U4892 ( .A(\CACHE[0][18] ), .B(\CACHE[1][18] ), .C(\CACHE[2][18] ), 
        .D(\CACHE[3][18] ), .S0(n3667), .S1(n3686), .Y(n3421) );
  MXI4X1 U4893 ( .A(\CACHE[4][18] ), .B(\CACHE[5][18] ), .C(\CACHE[6][18] ), 
        .D(\CACHE[7][18] ), .S0(n3666), .S1(n3705), .Y(n3422) );
  MXI4X1 U4894 ( .A(\CACHE[0][19] ), .B(\CACHE[1][19] ), .C(\CACHE[2][19] ), 
        .D(\CACHE[3][19] ), .S0(n3667), .S1(n3710), .Y(n3423) );
  MXI4X1 U4895 ( .A(\CACHE[4][19] ), .B(\CACHE[5][19] ), .C(\CACHE[6][19] ), 
        .D(\CACHE[7][19] ), .S0(n3667), .S1(n3695), .Y(n3424) );
  MXI4X1 U4896 ( .A(\CACHE[0][20] ), .B(\CACHE[1][20] ), .C(\CACHE[2][20] ), 
        .D(\CACHE[3][20] ), .S0(n3667), .S1(n3704), .Y(n3425) );
  MXI4X1 U4897 ( .A(\CACHE[4][20] ), .B(\CACHE[5][20] ), .C(\CACHE[6][20] ), 
        .D(\CACHE[7][20] ), .S0(n3667), .S1(n3699), .Y(n3426) );
  MXI4X1 U4898 ( .A(\CACHE[0][21] ), .B(\CACHE[1][21] ), .C(\CACHE[2][21] ), 
        .D(\CACHE[3][21] ), .S0(n3667), .S1(n3695), .Y(n3427) );
  MXI4X1 U4899 ( .A(\CACHE[4][21] ), .B(\CACHE[5][21] ), .C(\CACHE[6][21] ), 
        .D(\CACHE[7][21] ), .S0(n3667), .S1(n3700), .Y(n3428) );
  MXI4X1 U4900 ( .A(\CACHE[0][22] ), .B(\CACHE[1][22] ), .C(\CACHE[2][22] ), 
        .D(\CACHE[3][22] ), .S0(n3667), .S1(n3702), .Y(n3429) );
  MXI4X1 U4901 ( .A(\CACHE[4][22] ), .B(\CACHE[5][22] ), .C(\CACHE[6][22] ), 
        .D(\CACHE[7][22] ), .S0(n3667), .S1(n3697), .Y(n3430) );
  MXI4X1 U4902 ( .A(\CACHE[0][23] ), .B(\CACHE[1][23] ), .C(\CACHE[2][23] ), 
        .D(\CACHE[3][23] ), .S0(n3667), .S1(n3699), .Y(n3431) );
  MXI4X1 U4903 ( .A(\CACHE[4][23] ), .B(\CACHE[5][23] ), .C(\CACHE[6][23] ), 
        .D(\CACHE[7][23] ), .S0(n3667), .S1(n3699), .Y(n3432) );
  MXI4X1 U4904 ( .A(\CACHE[0][24] ), .B(\CACHE[1][24] ), .C(\CACHE[2][24] ), 
        .D(\CACHE[3][24] ), .S0(n3667), .S1(n3699), .Y(n3433) );
  MXI4X1 U4905 ( .A(\CACHE[4][24] ), .B(\CACHE[5][24] ), .C(\CACHE[6][24] ), 
        .D(\CACHE[7][24] ), .S0(n3667), .S1(n3699), .Y(n3434) );
  MXI4X1 U4906 ( .A(\CACHE[0][25] ), .B(\CACHE[1][25] ), .C(\CACHE[2][25] ), 
        .D(\CACHE[3][25] ), .S0(n3668), .S1(n3699), .Y(n3435) );
  MXI4X1 U4907 ( .A(\CACHE[4][25] ), .B(\CACHE[5][25] ), .C(\CACHE[6][25] ), 
        .D(\CACHE[7][25] ), .S0(n3668), .S1(n3699), .Y(n3436) );
  MXI4X1 U4908 ( .A(\CACHE[0][26] ), .B(\CACHE[1][26] ), .C(\CACHE[2][26] ), 
        .D(\CACHE[3][26] ), .S0(n3668), .S1(n3699), .Y(n3437) );
  MXI4X1 U4909 ( .A(\CACHE[4][26] ), .B(\CACHE[5][26] ), .C(\CACHE[6][26] ), 
        .D(\CACHE[7][26] ), .S0(n3668), .S1(n3699), .Y(n3438) );
  MXI4X1 U4910 ( .A(\CACHE[0][27] ), .B(\CACHE[1][27] ), .C(\CACHE[2][27] ), 
        .D(\CACHE[3][27] ), .S0(n3668), .S1(n3699), .Y(n3439) );
  MXI4X1 U4911 ( .A(\CACHE[4][27] ), .B(\CACHE[5][27] ), .C(\CACHE[6][27] ), 
        .D(\CACHE[7][27] ), .S0(n3668), .S1(n3699), .Y(n3440) );
  MXI4X1 U4912 ( .A(\CACHE[0][28] ), .B(\CACHE[1][28] ), .C(\CACHE[2][28] ), 
        .D(\CACHE[3][28] ), .S0(n3668), .S1(n3699), .Y(n3441) );
  MXI4X1 U4913 ( .A(\CACHE[4][28] ), .B(\CACHE[5][28] ), .C(\CACHE[6][28] ), 
        .D(\CACHE[7][28] ), .S0(n3668), .S1(n3699), .Y(n3442) );
  MXI4X1 U4914 ( .A(\CACHE[0][29] ), .B(\CACHE[1][29] ), .C(\CACHE[2][29] ), 
        .D(\CACHE[3][29] ), .S0(n3668), .S1(n3700), .Y(n3443) );
  MXI4X1 U4915 ( .A(\CACHE[4][29] ), .B(\CACHE[5][29] ), .C(\CACHE[6][29] ), 
        .D(\CACHE[7][29] ), .S0(n3668), .S1(n3700), .Y(n3444) );
  MXI4X1 U4916 ( .A(\CACHE[0][30] ), .B(\CACHE[1][30] ), .C(\CACHE[2][30] ), 
        .D(\CACHE[3][30] ), .S0(n3668), .S1(n3700), .Y(n3445) );
  MXI4X1 U4917 ( .A(\CACHE[4][30] ), .B(\CACHE[5][30] ), .C(\CACHE[6][30] ), 
        .D(\CACHE[7][30] ), .S0(n3668), .S1(n3700), .Y(n3446) );
  MXI4X1 U4918 ( .A(\CACHE[0][31] ), .B(\CACHE[1][31] ), .C(\CACHE[2][31] ), 
        .D(\CACHE[3][31] ), .S0(n3669), .S1(n3700), .Y(n3447) );
  MXI4X1 U4919 ( .A(\CACHE[4][31] ), .B(\CACHE[5][31] ), .C(\CACHE[6][31] ), 
        .D(\CACHE[7][31] ), .S0(n3668), .S1(n3700), .Y(n3448) );
  MXI4X1 U4920 ( .A(\CACHE[0][96] ), .B(\CACHE[1][96] ), .C(\CACHE[2][96] ), 
        .D(\CACHE[3][96] ), .S0(n3678), .S1(n3708), .Y(n3577) );
  MXI4X1 U4921 ( .A(\CACHE[4][96] ), .B(\CACHE[5][96] ), .C(\CACHE[6][96] ), 
        .D(\CACHE[7][96] ), .S0(n3677), .S1(n3708), .Y(n3578) );
  MXI4X1 U4922 ( .A(\CACHE[0][97] ), .B(\CACHE[1][97] ), .C(\CACHE[2][97] ), 
        .D(\CACHE[3][97] ), .S0(n3678), .S1(n3708), .Y(n3579) );
  MXI4X1 U4923 ( .A(\CACHE[4][97] ), .B(\CACHE[5][97] ), .C(\CACHE[6][97] ), 
        .D(\CACHE[7][97] ), .S0(n3678), .S1(n3708), .Y(n3580) );
  MXI4X1 U4924 ( .A(\CACHE[0][98] ), .B(\CACHE[1][98] ), .C(\CACHE[2][98] ), 
        .D(\CACHE[3][98] ), .S0(n3678), .S1(n3708), .Y(n3581) );
  MXI4X1 U4925 ( .A(\CACHE[4][98] ), .B(\CACHE[5][98] ), .C(\CACHE[6][98] ), 
        .D(\CACHE[7][98] ), .S0(n3678), .S1(n3708), .Y(n3582) );
  MXI4X1 U4926 ( .A(\CACHE[0][99] ), .B(\CACHE[1][99] ), .C(\CACHE[2][99] ), 
        .D(\CACHE[3][99] ), .S0(n3678), .S1(n3708), .Y(n3583) );
  MXI4X1 U4927 ( .A(\CACHE[4][99] ), .B(\CACHE[5][99] ), .C(\CACHE[6][99] ), 
        .D(\CACHE[7][99] ), .S0(n3678), .S1(n3708), .Y(n3584) );
  MXI4X1 U4928 ( .A(\CACHE[0][100] ), .B(\CACHE[1][100] ), .C(\CACHE[2][100] ), 
        .D(\CACHE[3][100] ), .S0(n3678), .S1(n3708), .Y(n3585) );
  MXI4X1 U4929 ( .A(\CACHE[4][100] ), .B(\CACHE[5][100] ), .C(\CACHE[6][100] ), 
        .D(\CACHE[7][100] ), .S0(n3678), .S1(n3708), .Y(n3586) );
  MXI4X1 U4930 ( .A(\CACHE[0][101] ), .B(\CACHE[1][101] ), .C(\CACHE[2][101] ), 
        .D(\CACHE[3][101] ), .S0(n3678), .S1(n3709), .Y(n3587) );
  MXI4X1 U4931 ( .A(\CACHE[4][101] ), .B(\CACHE[5][101] ), .C(\CACHE[6][101] ), 
        .D(\CACHE[7][101] ), .S0(n3678), .S1(n3709), .Y(n3588) );
  MXI4X1 U4932 ( .A(\CACHE[0][102] ), .B(\CACHE[1][102] ), .C(\CACHE[2][102] ), 
        .D(\CACHE[3][102] ), .S0(n3678), .S1(n3709), .Y(n3589) );
  MXI4X1 U4933 ( .A(\CACHE[4][102] ), .B(\CACHE[5][102] ), .C(\CACHE[6][102] ), 
        .D(\CACHE[7][102] ), .S0(n3678), .S1(n3709), .Y(n3590) );
  MXI4X1 U4934 ( .A(\CACHE[0][103] ), .B(\CACHE[1][103] ), .C(\CACHE[2][103] ), 
        .D(\CACHE[3][103] ), .S0(n3679), .S1(n3709), .Y(n3591) );
  MXI4X1 U4935 ( .A(\CACHE[4][103] ), .B(\CACHE[5][103] ), .C(\CACHE[6][103] ), 
        .D(\CACHE[7][103] ), .S0(n3679), .S1(n3709), .Y(n3592) );
  MXI4X1 U4936 ( .A(\CACHE[0][104] ), .B(\CACHE[1][104] ), .C(\CACHE[2][104] ), 
        .D(\CACHE[3][104] ), .S0(n3679), .S1(n3709), .Y(n3593) );
  MXI4X1 U4937 ( .A(\CACHE[4][104] ), .B(\CACHE[5][104] ), .C(\CACHE[6][104] ), 
        .D(\CACHE[7][104] ), .S0(n3679), .S1(n3709), .Y(n3594) );
  MXI4X1 U4938 ( .A(\CACHE[0][105] ), .B(\CACHE[1][105] ), .C(\CACHE[2][105] ), 
        .D(\CACHE[3][105] ), .S0(n3679), .S1(n3709), .Y(n3595) );
  MXI4X1 U4939 ( .A(\CACHE[4][105] ), .B(\CACHE[5][105] ), .C(\CACHE[6][105] ), 
        .D(\CACHE[7][105] ), .S0(n3679), .S1(n3709), .Y(n3596) );
  MXI4X1 U4940 ( .A(\CACHE[0][106] ), .B(\CACHE[1][106] ), .C(\CACHE[2][106] ), 
        .D(\CACHE[3][106] ), .S0(n3679), .S1(n3709), .Y(n3597) );
  MXI4X1 U4941 ( .A(\CACHE[4][106] ), .B(\CACHE[5][106] ), .C(\CACHE[6][106] ), 
        .D(\CACHE[7][106] ), .S0(n3679), .S1(n3709), .Y(n3598) );
  MXI4X1 U4942 ( .A(\CACHE[0][107] ), .B(\CACHE[1][107] ), .C(\CACHE[2][107] ), 
        .D(\CACHE[3][107] ), .S0(n3679), .S1(n3710), .Y(n3599) );
  MXI4X1 U4943 ( .A(\CACHE[4][107] ), .B(\CACHE[5][107] ), .C(\CACHE[6][107] ), 
        .D(\CACHE[7][107] ), .S0(n3679), .S1(n3710), .Y(n3600) );
  MXI4X1 U4944 ( .A(\CACHE[0][108] ), .B(\CACHE[1][108] ), .C(\CACHE[2][108] ), 
        .D(\CACHE[3][108] ), .S0(n3679), .S1(n3710), .Y(n3601) );
  MXI4X1 U4945 ( .A(\CACHE[4][108] ), .B(\CACHE[5][108] ), .C(\CACHE[6][108] ), 
        .D(\CACHE[7][108] ), .S0(n3679), .S1(n3710), .Y(n3602) );
  MXI4X1 U4946 ( .A(\CACHE[0][109] ), .B(\CACHE[1][109] ), .C(\CACHE[2][109] ), 
        .D(\CACHE[3][109] ), .S0(n3666), .S1(n3710), .Y(n3603) );
  MXI4X1 U4947 ( .A(\CACHE[4][109] ), .B(\CACHE[5][109] ), .C(\CACHE[6][109] ), 
        .D(\CACHE[7][109] ), .S0(n3679), .S1(n3710), .Y(n3604) );
  MXI4X1 U4948 ( .A(\CACHE[0][110] ), .B(\CACHE[1][110] ), .C(\CACHE[2][110] ), 
        .D(\CACHE[3][110] ), .S0(n3679), .S1(n3710), .Y(n3605) );
  MXI4X1 U4949 ( .A(\CACHE[4][110] ), .B(\CACHE[5][110] ), .C(\CACHE[6][110] ), 
        .D(\CACHE[7][110] ), .S0(n3667), .S1(n3710), .Y(n3606) );
  MXI4X1 U4950 ( .A(\CACHE[0][111] ), .B(\CACHE[1][111] ), .C(\CACHE[2][111] ), 
        .D(\CACHE[3][111] ), .S0(n3670), .S1(n3710), .Y(n3607) );
  MXI4X1 U4951 ( .A(\CACHE[4][111] ), .B(\CACHE[5][111] ), .C(\CACHE[6][111] ), 
        .D(\CACHE[7][111] ), .S0(n3677), .S1(n3710), .Y(n3608) );
  MXI4X1 U4952 ( .A(\CACHE[0][112] ), .B(\CACHE[1][112] ), .C(\CACHE[2][112] ), 
        .D(\CACHE[3][112] ), .S0(n3669), .S1(n3710), .Y(n3609) );
  MXI4X1 U4953 ( .A(\CACHE[4][112] ), .B(\CACHE[5][112] ), .C(\CACHE[6][112] ), 
        .D(\CACHE[7][112] ), .S0(n3672), .S1(n3710), .Y(n3610) );
  MXI4X1 U4954 ( .A(\CACHE[0][113] ), .B(\CACHE[1][113] ), .C(\CACHE[2][113] ), 
        .D(\CACHE[3][113] ), .S0(n3674), .S1(n3710), .Y(n3611) );
  MXI4X1 U4955 ( .A(\CACHE[4][113] ), .B(\CACHE[5][113] ), .C(\CACHE[6][113] ), 
        .D(\CACHE[7][113] ), .S0(n3679), .S1(n3699), .Y(n3612) );
  MXI4X1 U4956 ( .A(\CACHE[0][114] ), .B(\CACHE[1][114] ), .C(\CACHE[2][114] ), 
        .D(\CACHE[3][114] ), .S0(n3676), .S1(n3700), .Y(n3613) );
  MXI4X1 U4957 ( .A(\CACHE[4][114] ), .B(\CACHE[5][114] ), .C(\CACHE[6][114] ), 
        .D(\CACHE[7][114] ), .S0(n3666), .S1(n3700), .Y(n3614) );
  MXI4X1 U4958 ( .A(\CACHE[0][115] ), .B(\CACHE[1][115] ), .C(\CACHE[2][115] ), 
        .D(\CACHE[3][115] ), .S0(n3675), .S1(n3699), .Y(n3615) );
  MXI4X1 U4959 ( .A(\CACHE[4][115] ), .B(\CACHE[5][115] ), .C(\CACHE[6][115] ), 
        .D(\CACHE[7][115] ), .S0(n3678), .S1(n3699), .Y(n3616) );
  MXI4X1 U4960 ( .A(\CACHE[0][116] ), .B(\CACHE[1][116] ), .C(\CACHE[2][116] ), 
        .D(\CACHE[3][116] ), .S0(n3680), .S1(n3710), .Y(n3617) );
  MXI4X1 U4961 ( .A(\CACHE[4][116] ), .B(\CACHE[5][116] ), .C(\CACHE[6][116] ), 
        .D(\CACHE[7][116] ), .S0(n3680), .S1(n3710), .Y(n3618) );
  MXI4X1 U4962 ( .A(\CACHE[0][117] ), .B(\CACHE[1][117] ), .C(\CACHE[2][117] ), 
        .D(\CACHE[3][117] ), .S0(n3680), .S1(n3700), .Y(n3619) );
  MXI4X1 U4963 ( .A(\CACHE[4][117] ), .B(\CACHE[5][117] ), .C(\CACHE[6][117] ), 
        .D(\CACHE[7][117] ), .S0(n3680), .S1(n3700), .Y(n3620) );
  MXI4X1 U4964 ( .A(\CACHE[0][118] ), .B(\CACHE[1][118] ), .C(\CACHE[2][118] ), 
        .D(\CACHE[3][118] ), .S0(n3680), .S1(n3699), .Y(n3621) );
  MXI4X1 U4965 ( .A(\CACHE[4][118] ), .B(\CACHE[5][118] ), .C(\CACHE[6][118] ), 
        .D(\CACHE[7][118] ), .S0(n3680), .S1(n3710), .Y(n3622) );
  INVX3 U4966 ( .A(proc_reset), .Y(n4142) );
endmodule

