
module IFID ( IF_Flush, clk, IFIDWrite, PC_plus4, PC_plus4Reg, Inst, InstReg, 
        stall_bothzero );
  input [31:0] PC_plus4;
  output [31:0] PC_plus4Reg;
  input [31:0] Inst;
  output [31:0] InstReg;
  input IF_Flush, clk, IFIDWrite, stall_bothzero;
  wire   N3, n1, n3, n5, n7, n9, n11, n13;
  wire   [31:0] IF_pcplus4;
  wire   [31:0] IF_Inst;

  EDFFX1 \PC_plus4Reg_reg[1]  ( .D(IF_pcplus4[1]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[1]) );
  EDFFX1 \PC_plus4Reg_reg[0]  ( .D(IF_pcplus4[0]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[0]) );
  EDFFX1 \PC_plus4Reg_reg[27]  ( .D(IF_pcplus4[27]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[27]) );
  EDFFX1 \PC_plus4Reg_reg[26]  ( .D(IF_pcplus4[26]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[26]) );
  EDFFX1 \PC_plus4Reg_reg[25]  ( .D(IF_pcplus4[25]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[25]) );
  EDFFX1 \PC_plus4Reg_reg[24]  ( .D(IF_pcplus4[24]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[24]) );
  EDFFX1 \PC_plus4Reg_reg[23]  ( .D(IF_pcplus4[23]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[23]) );
  EDFFX1 \PC_plus4Reg_reg[22]  ( .D(IF_pcplus4[22]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[22]) );
  EDFFX1 \PC_plus4Reg_reg[21]  ( .D(IF_pcplus4[21]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[21]) );
  EDFFX1 \PC_plus4Reg_reg[20]  ( .D(IF_pcplus4[20]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[20]) );
  EDFFX1 \PC_plus4Reg_reg[19]  ( .D(IF_pcplus4[19]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[19]) );
  EDFFX1 \PC_plus4Reg_reg[18]  ( .D(IF_pcplus4[18]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[18]) );
  EDFFX1 \PC_plus4Reg_reg[17]  ( .D(IF_pcplus4[17]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[17]) );
  EDFFX1 \PC_plus4Reg_reg[16]  ( .D(IF_pcplus4[16]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[16]) );
  EDFFX1 \PC_plus4Reg_reg[15]  ( .D(IF_pcplus4[15]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[15]) );
  EDFFX1 \PC_plus4Reg_reg[14]  ( .D(IF_pcplus4[14]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[14]) );
  EDFFX1 \PC_plus4Reg_reg[13]  ( .D(IF_pcplus4[13]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[13]) );
  EDFFX1 \PC_plus4Reg_reg[12]  ( .D(IF_pcplus4[12]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[12]) );
  EDFFX1 \PC_plus4Reg_reg[11]  ( .D(IF_pcplus4[11]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[11]) );
  EDFFX1 \PC_plus4Reg_reg[10]  ( .D(IF_pcplus4[10]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[10]) );
  EDFFX1 \PC_plus4Reg_reg[9]  ( .D(IF_pcplus4[9]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[9]) );
  EDFFX1 \PC_plus4Reg_reg[8]  ( .D(IF_pcplus4[8]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[8]) );
  EDFFX1 \PC_plus4Reg_reg[7]  ( .D(IF_pcplus4[7]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[7]) );
  EDFFX1 \PC_plus4Reg_reg[6]  ( .D(IF_pcplus4[6]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[6]) );
  EDFFX1 \PC_plus4Reg_reg[5]  ( .D(IF_pcplus4[5]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[5]) );
  EDFFX1 \PC_plus4Reg_reg[4]  ( .D(IF_pcplus4[4]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[4]) );
  EDFFX1 \PC_plus4Reg_reg[3]  ( .D(IF_pcplus4[3]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[3]) );
  EDFFX1 \PC_plus4Reg_reg[31]  ( .D(IF_pcplus4[31]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[31]) );
  EDFFX1 \PC_plus4Reg_reg[30]  ( .D(IF_pcplus4[30]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[30]) );
  EDFFX1 \PC_plus4Reg_reg[29]  ( .D(IF_pcplus4[29]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[29]) );
  EDFFX1 \PC_plus4Reg_reg[28]  ( .D(IF_pcplus4[28]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[28]) );
  EDFFX1 \InstReg_reg[27]  ( .D(IF_Inst[27]), .E(N3), .CK(clk), .Q(InstReg[27]) );
  EDFFX1 \PC_plus4Reg_reg[2]  ( .D(IF_pcplus4[2]), .E(N3), .CK(clk), .Q(
        PC_plus4Reg[2]) );
  EDFFX1 \InstReg_reg[30]  ( .D(IF_Inst[30]), .E(N3), .CK(clk), .Q(InstReg[30]) );
  EDFFX1 \InstReg_reg[28]  ( .D(IF_Inst[28]), .E(N3), .CK(clk), .Q(InstReg[28]) );
  EDFFX1 \InstReg_reg[0]  ( .D(IF_Inst[0]), .E(N3), .CK(clk), .Q(InstReg[0])
         );
  EDFFX1 \InstReg_reg[10]  ( .D(IF_Inst[10]), .E(N3), .CK(clk), .Q(InstReg[10]) );
  EDFFX1 \InstReg_reg[9]  ( .D(IF_Inst[9]), .E(N3), .CK(clk), .Q(InstReg[9])
         );
  EDFFX1 \InstReg_reg[8]  ( .D(IF_Inst[8]), .E(N3), .CK(clk), .Q(InstReg[8])
         );
  EDFFX1 \InstReg_reg[7]  ( .D(IF_Inst[7]), .E(N3), .CK(clk), .Q(InstReg[7])
         );
  EDFFX1 \InstReg_reg[6]  ( .D(IF_Inst[6]), .E(N3), .CK(clk), .Q(InstReg[6])
         );
  EDFFX1 \InstReg_reg[5]  ( .D(IF_Inst[5]), .E(N3), .CK(clk), .Q(InstReg[5])
         );
  EDFFX1 \InstReg_reg[4]  ( .D(IF_Inst[4]), .E(N3), .CK(clk), .Q(InstReg[4])
         );
  EDFFX1 \InstReg_reg[3]  ( .D(IF_Inst[3]), .E(N3), .CK(clk), .Q(InstReg[3])
         );
  EDFFX1 \InstReg_reg[2]  ( .D(IF_Inst[2]), .E(N3), .CK(clk), .Q(InstReg[2])
         );
  EDFFX1 \InstReg_reg[1]  ( .D(IF_Inst[1]), .E(N3), .CK(clk), .Q(InstReg[1])
         );
  EDFFX1 \InstReg_reg[26]  ( .D(IF_Inst[26]), .E(N3), .CK(clk), .Q(InstReg[26]) );
  EDFFX1 \InstReg_reg[31]  ( .D(IF_Inst[31]), .E(N3), .CK(clk), .Q(InstReg[31]) );
  EDFFX1 \InstReg_reg[11]  ( .D(IF_Inst[11]), .E(N3), .CK(clk), .Q(InstReg[11]) );
  EDFFX1 \InstReg_reg[12]  ( .D(IF_Inst[12]), .E(N3), .CK(clk), .Q(InstReg[12]) );
  EDFFX1 \InstReg_reg[13]  ( .D(IF_Inst[13]), .E(N3), .CK(clk), .Q(InstReg[13]) );
  EDFFX1 \InstReg_reg[14]  ( .D(IF_Inst[14]), .E(N3), .CK(clk), .Q(InstReg[14]) );
  EDFFX1 \InstReg_reg[22]  ( .D(IF_Inst[22]), .E(N3), .CK(clk), .Q(InstReg[22]) );
  EDFFX1 \InstReg_reg[17]  ( .D(IF_Inst[17]), .E(N3), .CK(clk), .Q(InstReg[17]) );
  EDFFX2 \InstReg_reg[29]  ( .D(IF_Inst[29]), .E(N3), .CK(clk), .Q(InstReg[29]) );
  EDFFX1 \InstReg_reg[21]  ( .D(IF_Inst[21]), .E(N3), .CK(clk), .Q(InstReg[21]) );
  EDFFX1 \InstReg_reg[16]  ( .D(IF_Inst[16]), .E(N3), .CK(clk), .Q(InstReg[16]) );
  EDFFX1 \InstReg_reg[24]  ( .D(IF_Inst[24]), .E(N3), .CK(clk), .QN(n13) );
  EDFFX1 \InstReg_reg[19]  ( .D(IF_Inst[19]), .E(N3), .CK(clk), .QN(n11) );
  EDFFX1 \InstReg_reg[23]  ( .D(IF_Inst[23]), .E(N3), .CK(clk), .QN(n9) );
  EDFFX1 \InstReg_reg[18]  ( .D(IF_Inst[18]), .E(N3), .CK(clk), .QN(n7) );
  EDFFX1 \InstReg_reg[25]  ( .D(IF_Inst[25]), .E(N3), .CK(clk), .QN(n5) );
  EDFFX1 \InstReg_reg[20]  ( .D(IF_Inst[20]), .E(N3), .CK(clk), .QN(n3) );
  EDFFX1 \InstReg_reg[15]  ( .D(IF_Inst[15]), .E(N3), .CK(clk), .QN(n1) );
  CLKAND2X12 U2 ( .A(stall_bothzero), .B(IFIDWrite), .Y(N3) );
  INVX6 U3 ( .A(n1), .Y(InstReg[15]) );
  INVX6 U4 ( .A(n3), .Y(InstReg[20]) );
  INVX8 U5 ( .A(n5), .Y(InstReg[25]) );
  INVX12 U6 ( .A(n7), .Y(InstReg[18]) );
  INVX12 U7 ( .A(n9), .Y(InstReg[23]) );
  INVX16 U8 ( .A(n11), .Y(InstReg[19]) );
  INVX16 U9 ( .A(n13), .Y(InstReg[24]) );
  NOR2BXL U10 ( .AN(Inst[15]), .B(IF_Flush), .Y(IF_Inst[15]) );
  NOR2BXL U11 ( .AN(Inst[18]), .B(IF_Flush), .Y(IF_Inst[18]) );
  NOR2BXL U12 ( .AN(Inst[19]), .B(IF_Flush), .Y(IF_Inst[19]) );
  NOR2BXL U13 ( .AN(Inst[20]), .B(IF_Flush), .Y(IF_Inst[20]) );
  NOR2BXL U14 ( .AN(Inst[23]), .B(IF_Flush), .Y(IF_Inst[23]) );
  NOR2BXL U15 ( .AN(Inst[24]), .B(IF_Flush), .Y(IF_Inst[24]) );
  NOR2BXL U16 ( .AN(Inst[25]), .B(IF_Flush), .Y(IF_Inst[25]) );
  NOR2BXL U17 ( .AN(Inst[29]), .B(IF_Flush), .Y(IF_Inst[29]) );
  NOR2BXL U18 ( .AN(PC_plus4[0]), .B(IF_Flush), .Y(IF_pcplus4[0]) );
  NOR2BXL U19 ( .AN(PC_plus4[1]), .B(IF_Flush), .Y(IF_pcplus4[1]) );
  NOR2BXL U20 ( .AN(PC_plus4[2]), .B(IF_Flush), .Y(IF_pcplus4[2]) );
  NOR2BXL U21 ( .AN(PC_plus4[3]), .B(IF_Flush), .Y(IF_pcplus4[3]) );
  NOR2BXL U22 ( .AN(PC_plus4[4]), .B(IF_Flush), .Y(IF_pcplus4[4]) );
  NOR2BXL U23 ( .AN(PC_plus4[5]), .B(IF_Flush), .Y(IF_pcplus4[5]) );
  NOR2BXL U24 ( .AN(PC_plus4[6]), .B(IF_Flush), .Y(IF_pcplus4[6]) );
  NOR2BXL U25 ( .AN(PC_plus4[7]), .B(IF_Flush), .Y(IF_pcplus4[7]) );
  NOR2BXL U26 ( .AN(PC_plus4[8]), .B(IF_Flush), .Y(IF_pcplus4[8]) );
  NOR2BXL U27 ( .AN(PC_plus4[9]), .B(IF_Flush), .Y(IF_pcplus4[9]) );
  NOR2BXL U28 ( .AN(PC_plus4[10]), .B(IF_Flush), .Y(IF_pcplus4[10]) );
  NOR2BXL U29 ( .AN(PC_plus4[11]), .B(IF_Flush), .Y(IF_pcplus4[11]) );
  NOR2BXL U30 ( .AN(PC_plus4[12]), .B(IF_Flush), .Y(IF_pcplus4[12]) );
  NOR2BXL U31 ( .AN(PC_plus4[13]), .B(IF_Flush), .Y(IF_pcplus4[13]) );
  NOR2BXL U32 ( .AN(PC_plus4[14]), .B(IF_Flush), .Y(IF_pcplus4[14]) );
  NOR2BXL U33 ( .AN(PC_plus4[15]), .B(IF_Flush), .Y(IF_pcplus4[15]) );
  NOR2BXL U34 ( .AN(PC_plus4[16]), .B(IF_Flush), .Y(IF_pcplus4[16]) );
  NOR2BXL U35 ( .AN(PC_plus4[17]), .B(IF_Flush), .Y(IF_pcplus4[17]) );
  NOR2BXL U36 ( .AN(PC_plus4[18]), .B(IF_Flush), .Y(IF_pcplus4[18]) );
  NOR2BXL U37 ( .AN(PC_plus4[19]), .B(IF_Flush), .Y(IF_pcplus4[19]) );
  NOR2BXL U38 ( .AN(PC_plus4[20]), .B(IF_Flush), .Y(IF_pcplus4[20]) );
  NOR2BXL U39 ( .AN(PC_plus4[21]), .B(IF_Flush), .Y(IF_pcplus4[21]) );
  NOR2BXL U40 ( .AN(PC_plus4[22]), .B(IF_Flush), .Y(IF_pcplus4[22]) );
  NOR2BXL U41 ( .AN(PC_plus4[23]), .B(IF_Flush), .Y(IF_pcplus4[23]) );
  NOR2BXL U42 ( .AN(PC_plus4[24]), .B(IF_Flush), .Y(IF_pcplus4[24]) );
  NOR2BXL U43 ( .AN(PC_plus4[25]), .B(IF_Flush), .Y(IF_pcplus4[25]) );
  NOR2BXL U44 ( .AN(PC_plus4[26]), .B(IF_Flush), .Y(IF_pcplus4[26]) );
  NOR2BXL U45 ( .AN(PC_plus4[27]), .B(IF_Flush), .Y(IF_pcplus4[27]) );
  NOR2BXL U46 ( .AN(PC_plus4[28]), .B(IF_Flush), .Y(IF_pcplus4[28]) );
  NOR2BXL U47 ( .AN(PC_plus4[29]), .B(IF_Flush), .Y(IF_pcplus4[29]) );
  NOR2BXL U48 ( .AN(PC_plus4[30]), .B(IF_Flush), .Y(IF_pcplus4[30]) );
  NOR2BXL U49 ( .AN(PC_plus4[31]), .B(IF_Flush), .Y(IF_pcplus4[31]) );
  NOR2BXL U50 ( .AN(Inst[0]), .B(IF_Flush), .Y(IF_Inst[0]) );
  NOR2BXL U51 ( .AN(Inst[1]), .B(IF_Flush), .Y(IF_Inst[1]) );
  NOR2BXL U52 ( .AN(Inst[2]), .B(IF_Flush), .Y(IF_Inst[2]) );
  NOR2BXL U53 ( .AN(Inst[3]), .B(IF_Flush), .Y(IF_Inst[3]) );
  NOR2BXL U54 ( .AN(Inst[4]), .B(IF_Flush), .Y(IF_Inst[4]) );
  NOR2BXL U55 ( .AN(Inst[5]), .B(IF_Flush), .Y(IF_Inst[5]) );
  NOR2BXL U56 ( .AN(Inst[6]), .B(IF_Flush), .Y(IF_Inst[6]) );
  NOR2BXL U57 ( .AN(Inst[7]), .B(IF_Flush), .Y(IF_Inst[7]) );
  NOR2BXL U58 ( .AN(Inst[8]), .B(IF_Flush), .Y(IF_Inst[8]) );
  NOR2BXL U59 ( .AN(Inst[9]), .B(IF_Flush), .Y(IF_Inst[9]) );
  NOR2BXL U60 ( .AN(Inst[10]), .B(IF_Flush), .Y(IF_Inst[10]) );
  NOR2BXL U61 ( .AN(Inst[11]), .B(IF_Flush), .Y(IF_Inst[11]) );
  NOR2BXL U62 ( .AN(Inst[12]), .B(IF_Flush), .Y(IF_Inst[12]) );
  NOR2BXL U63 ( .AN(Inst[13]), .B(IF_Flush), .Y(IF_Inst[13]) );
  NOR2BXL U64 ( .AN(Inst[14]), .B(IF_Flush), .Y(IF_Inst[14]) );
  NOR2BXL U65 ( .AN(Inst[16]), .B(IF_Flush), .Y(IF_Inst[16]) );
  NOR2BXL U66 ( .AN(Inst[17]), .B(IF_Flush), .Y(IF_Inst[17]) );
  NOR2BXL U67 ( .AN(Inst[21]), .B(IF_Flush), .Y(IF_Inst[21]) );
  NOR2BXL U68 ( .AN(Inst[22]), .B(IF_Flush), .Y(IF_Inst[22]) );
  NOR2BXL U69 ( .AN(Inst[26]), .B(IF_Flush), .Y(IF_Inst[26]) );
  NOR2BXL U70 ( .AN(Inst[27]), .B(IF_Flush), .Y(IF_Inst[27]) );
  NOR2BXL U71 ( .AN(Inst[28]), .B(IF_Flush), .Y(IF_Inst[28]) );
  NOR2BXL U72 ( .AN(Inst[30]), .B(IF_Flush), .Y(IF_Inst[30]) );
  NOR2BXL U73 ( .AN(Inst[31]), .B(IF_Flush), .Y(IF_Inst[31]) );
endmodule


module Hazard_detection ( IDRegRS, IDRegRt, EXRegRt, EXMemRead, PCWrite, 
        IFIDWrite, HazMux );
  input [4:0] IDRegRS;
  input [4:0] IDRegRt;
  input [4:0] EXRegRt;
  input EXMemRead;
  output PCWrite, IFIDWrite, HazMux;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  XNOR2XL U1 ( .A(EXRegRt[3]), .B(IDRegRt[3]), .Y(n13) );
  XNOR2XL U2 ( .A(EXRegRt[3]), .B(IDRegRS[3]), .Y(n10) );
  XOR2XL U3 ( .A(IDRegRS[2]), .B(EXRegRt[2]), .Y(n8) );
  XOR2XL U4 ( .A(IDRegRt[2]), .B(EXRegRt[2]), .Y(n5) );
  XOR2XL U5 ( .A(IDRegRt[4]), .B(EXRegRt[4]), .Y(n6) );
  XOR2XL U6 ( .A(IDRegRS[4]), .B(EXRegRt[4]), .Y(n9) );
  BUFX2 U7 ( .A(IFIDWrite), .Y(PCWrite) );
  BUFX2 U8 ( .A(IFIDWrite), .Y(HazMux) );
  NAND2X1 U9 ( .A(EXMemRead), .B(n3), .Y(IFIDWrite) );
  OAI33X1 U10 ( .A0(n4), .A1(n5), .A2(n6), .B0(n7), .B1(n8), .B2(n9), .Y(n3)
         );
  NAND3X1 U11 ( .A(n10), .B(n11), .C(n12), .Y(n7) );
  XNOR2X1 U12 ( .A(EXRegRt[0]), .B(IDRegRS[0]), .Y(n12) );
  XNOR2X1 U13 ( .A(EXRegRt[1]), .B(IDRegRS[1]), .Y(n11) );
  NAND3X1 U14 ( .A(n13), .B(n14), .C(n15), .Y(n4) );
  XNOR2X1 U15 ( .A(EXRegRt[0]), .B(IDRegRt[0]), .Y(n15) );
  XNOR2X1 U16 ( .A(EXRegRt[1]), .B(IDRegRt[1]), .Y(n14) );
endmodule


module control ( opcode, rst_n, Rs, Rt, Rd, RegDST, MemtoReg, Jump, Branch, 
        MemRead, MemWrite, ALUSrc, RegWrite, ALUOp );
  input [5:0] opcode;
  input [4:0] Rs;
  input [4:0] Rt;
  input [4:0] Rd;
  output [1:0] RegDST;
  output [1:0] MemtoReg;
  output [1:0] Jump;
  output [2:0] ALUOp;
  input rst_n;
  output Branch, MemRead, MemWrite, ALUSrc, RegWrite;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37;

  NOR4X2 U3 ( .A(n2), .B(opcode[0]), .C(opcode[4]), .D(opcode[5]), .Y(n18) );
  OAI31X1 U4 ( .A0(n14), .A1(opcode[3]), .A2(opcode[2]), .B0(n10), .Y(Jump[1])
         );
  NAND2BXL U5 ( .AN(n23), .B(n24), .Y(n6) );
  NAND4XL U6 ( .A(n18), .B(n7), .C(n22), .D(n12), .Y(n11) );
  NAND3XL U7 ( .A(n22), .B(n21), .C(n18), .Y(n31) );
  AOI22XL U8 ( .A0(n15), .A1(n16), .B0(n17), .B1(n18), .Y(n14) );
  NOR4XL U9 ( .A(Rs[1]), .B(Rs[0]), .C(Rs[2]), .D(n32), .Y(n23) );
  OR2XL U10 ( .A(Rs[4]), .B(Rs[3]), .Y(n32) );
  NAND4XL U11 ( .A(opcode[2]), .B(n18), .C(n22), .D(n12), .Y(n19) );
  NOR3XL U12 ( .A(Rt[2]), .B(Rt[4]), .C(Rt[3]), .Y(n36) );
  NAND2XL U13 ( .A(opcode[3]), .B(n18), .Y(n26) );
  NOR3XL U14 ( .A(Rd[2]), .B(Rd[4]), .C(Rd[3]), .Y(n34) );
  CLKINVX1 U15 ( .A(rst_n), .Y(n2) );
  BUFX2 U16 ( .A(RegDST[1]), .Y(MemtoReg[1]) );
  OAI221XL U17 ( .A0(opcode[3]), .A1(n3), .B0(opcode[5]), .B1(n4), .C0(n5), 
        .Y(RegWrite) );
  AOI31X1 U18 ( .A0(n6), .A1(n7), .A2(n8), .B0(n9), .Y(n5) );
  OAI31XL U19 ( .A0(n3), .A1(opcode[5]), .A2(opcode[3]), .B0(n10), .Y(
        RegDST[1]) );
  CLKINVX1 U20 ( .A(n11), .Y(RegDST[0]) );
  NOR2X1 U21 ( .A(n12), .B(n13), .Y(MemWrite) );
  NOR2X1 U22 ( .A(opcode[3]), .B(n13), .Y(MemRead) );
  CLKINVX1 U23 ( .A(n6), .Y(n17) );
  OAI211X1 U24 ( .A0(n6), .A1(n11), .B0(n19), .C0(n10), .Y(Jump[0]) );
  NAND4X1 U25 ( .A(n20), .B(opcode[0]), .C(n21), .D(n16), .Y(n10) );
  CLKINVX1 U26 ( .A(n19), .Y(Branch) );
  NAND3X1 U27 ( .A(n25), .B(n13), .C(n26), .Y(ALUSrc) );
  CLKINVX1 U28 ( .A(MemtoReg[0]), .Y(n13) );
  NOR2X1 U29 ( .A(n16), .B(n3), .Y(MemtoReg[0]) );
  NAND3X1 U30 ( .A(n15), .B(n21), .C(opcode[0]), .Y(n3) );
  NOR3X1 U31 ( .A(n2), .B(opcode[4]), .C(n22), .Y(n15) );
  CLKINVX1 U32 ( .A(opcode[5]), .Y(n16) );
  OAI211X1 U33 ( .A0(n7), .A1(n27), .B0(n28), .C0(n25), .Y(ALUOp[2]) );
  CLKINVX1 U34 ( .A(n29), .Y(n25) );
  NAND2X1 U35 ( .A(n8), .B(n12), .Y(n27) );
  OAI221XL U36 ( .A0(n30), .A1(n31), .B0(opcode[2]), .B1(n26), .C0(n28), .Y(
        ALUOp[1]) );
  CLKINVX1 U37 ( .A(n7), .Y(n30) );
  NAND2X1 U38 ( .A(n24), .B(n23), .Y(n7) );
  AND4X1 U39 ( .A(n33), .B(n34), .C(n35), .D(n36), .Y(n24) );
  NOR2X1 U40 ( .A(Rt[1]), .B(Rt[0]), .Y(n35) );
  NOR2X1 U41 ( .A(Rd[1]), .B(Rd[0]), .Y(n33) );
  OAI211X1 U42 ( .A0(n21), .A1(n28), .B0(n19), .C0(n37), .Y(ALUOp[0]) );
  AOI22X1 U43 ( .A0(n29), .A1(opcode[0]), .B0(n8), .B1(opcode[3]), .Y(n37) );
  CLKINVX1 U44 ( .A(n31), .Y(n8) );
  NOR3X1 U45 ( .A(n4), .B(opcode[5]), .C(n21), .Y(n29) );
  CLKINVX1 U46 ( .A(n20), .Y(n4) );
  NOR4X1 U47 ( .A(n12), .B(n2), .C(opcode[1]), .D(opcode[4]), .Y(n20) );
  CLKINVX1 U48 ( .A(opcode[3]), .Y(n12) );
  CLKINVX1 U49 ( .A(opcode[1]), .Y(n22) );
  NAND2X1 U50 ( .A(n9), .B(opcode[1]), .Y(n28) );
  CLKINVX1 U51 ( .A(n26), .Y(n9) );
  CLKINVX1 U52 ( .A(opcode[2]), .Y(n21) );
endmodule


module beq_foward ( RegWrite, instruction31_26, instruction25_21, 
        instruction20_16, EX_Rd, Foward_C, Foward_D );
  input [5:0] instruction31_26;
  input [4:0] instruction25_21;
  input [4:0] instruction20_16;
  input [4:0] EX_Rd;
  input RegWrite;
  output Foward_C, Foward_D;
  wire   n18, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17;

  INVX6 U1 ( .A(n9), .Y(Foward_C) );
  NAND4XL U2 ( .A(n10), .B(n8), .C(n11), .D(n12), .Y(n9) );
  CLKBUFX6 U3 ( .A(n18), .Y(Foward_D) );
  XNOR2XL U4 ( .A(EX_Rd[3]), .B(instruction20_16[3]), .Y(n7) );
  XOR2XL U5 ( .A(instruction20_16[2]), .B(EX_Rd[2]), .Y(n5) );
  XOR2XL U6 ( .A(instruction20_16[4]), .B(EX_Rd[4]), .Y(n3) );
  XOR2XL U7 ( .A(instruction25_21[3]), .B(EX_Rd[3]), .Y(n13) );
  XOR2XL U8 ( .A(instruction25_21[2]), .B(EX_Rd[2]), .Y(n15) );
  XOR2XL U9 ( .A(instruction25_21[4]), .B(EX_Rd[4]), .Y(n14) );
  NOR4X1 U10 ( .A(n2), .B(n3), .C(n4), .D(n5), .Y(n18) );
  XOR2X1 U11 ( .A(instruction20_16[1]), .B(EX_Rd[1]), .Y(n4) );
  NAND4X1 U12 ( .A(n6), .B(n7), .C(n8), .D(n9), .Y(n2) );
  XNOR2X1 U13 ( .A(EX_Rd[0]), .B(instruction20_16[0]), .Y(n6) );
  NOR3X1 U14 ( .A(n13), .B(n14), .C(n15), .Y(n12) );
  XNOR2X1 U15 ( .A(EX_Rd[0]), .B(instruction25_21[0]), .Y(n11) );
  AND4X1 U16 ( .A(n16), .B(RegWrite), .C(instruction31_26[2]), .D(n17), .Y(n8)
         );
  NOR4X1 U17 ( .A(instruction31_26[5]), .B(instruction31_26[4]), .C(
        instruction31_26[3]), .D(instruction31_26[1]), .Y(n17) );
  CLKINVX1 U18 ( .A(instruction31_26[0]), .Y(n16) );
  XNOR2X1 U19 ( .A(EX_Rd[1]), .B(instruction25_21[1]), .Y(n10) );
endmodule


module IDEX ( clk, WB, M, EX, RegRs, RegRt, RegRd, data1, data2, sign_extend, 
        PC_plus4Reg, WB_reg, M_reg, EX_reg, RegRs_reg, RegRt_reg, RegRd_reg, 
        data1_reg, data2_reg, EX_pcplus4, sign_extend_reg, stall_bothzero );
  input [2:0] WB;
  input [2:0] M;
  input [5:0] EX;
  input [4:0] RegRs;
  input [4:0] RegRt;
  input [4:0] RegRd;
  input [31:0] data1;
  input [31:0] data2;
  input [31:0] sign_extend;
  input [31:0] PC_plus4Reg;
  output [2:0] WB_reg;
  output [2:0] M_reg;
  output [5:0] EX_reg;
  output [4:0] RegRs_reg;
  output [4:0] RegRt_reg;
  output [4:0] RegRd_reg;
  output [31:0] data1_reg;
  output [31:0] data2_reg;
  output [31:0] EX_pcplus4;
  output [31:0] sign_extend_reg;
  input clk, stall_bothzero;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  EDFFX1 \EX_reg_reg[0]  ( .D(EX[0]), .E(n9), .CK(clk), .Q(EX_reg[0]) );
  EDFFX1 \EX_reg_reg[4]  ( .D(EX[4]), .E(n10), .CK(clk), .Q(EX_reg[4]) );
  EDFFX1 \EX_reg_reg[2]  ( .D(EX[2]), .E(n9), .CK(clk), .Q(EX_reg[2]) );
  EDFFX1 \EX_reg_reg[1]  ( .D(EX[1]), .E(n9), .CK(clk), .Q(EX_reg[1]) );
  EDFFX1 \data1_reg_reg[31]  ( .D(data1[31]), .E(n3), .CK(clk), .Q(
        data1_reg[31]) );
  EDFFX1 \data1_reg_reg[30]  ( .D(data1[30]), .E(n3), .CK(clk), .Q(
        data1_reg[30]) );
  EDFFX1 \data1_reg_reg[29]  ( .D(data1[29]), .E(n3), .CK(clk), .Q(
        data1_reg[29]) );
  EDFFX1 \data1_reg_reg[28]  ( .D(data1[28]), .E(n3), .CK(clk), .Q(
        data1_reg[28]) );
  EDFFX1 \data1_reg_reg[27]  ( .D(data1[27]), .E(n4), .CK(clk), .Q(
        data1_reg[27]) );
  EDFFX1 \data1_reg_reg[26]  ( .D(data1[26]), .E(n4), .CK(clk), .Q(
        data1_reg[26]) );
  EDFFX1 \data1_reg_reg[25]  ( .D(data1[25]), .E(n4), .CK(clk), .Q(
        data1_reg[25]) );
  EDFFX1 \data1_reg_reg[24]  ( .D(data1[24]), .E(n4), .CK(clk), .Q(
        data1_reg[24]) );
  EDFFX1 \data1_reg_reg[23]  ( .D(data1[23]), .E(n5), .CK(clk), .Q(
        data1_reg[23]) );
  EDFFX1 \data1_reg_reg[22]  ( .D(data1[22]), .E(n5), .CK(clk), .Q(
        data1_reg[22]) );
  EDFFX1 \data1_reg_reg[21]  ( .D(data1[21]), .E(n5), .CK(clk), .Q(
        data1_reg[21]) );
  EDFFX1 \data1_reg_reg[20]  ( .D(data1[20]), .E(n5), .CK(clk), .Q(
        data1_reg[20]) );
  EDFFX1 \data1_reg_reg[19]  ( .D(data1[19]), .E(n5), .CK(clk), .Q(
        data1_reg[19]) );
  EDFFX1 \data1_reg_reg[18]  ( .D(data1[18]), .E(n14), .CK(clk), .Q(
        data1_reg[18]) );
  EDFFX1 \data1_reg_reg[17]  ( .D(data1[17]), .E(n6), .CK(clk), .Q(
        data1_reg[17]) );
  EDFFX1 \data1_reg_reg[16]  ( .D(data1[16]), .E(n6), .CK(clk), .Q(
        data1_reg[16]) );
  EDFFX1 \data1_reg_reg[15]  ( .D(data1[15]), .E(n6), .CK(clk), .Q(
        data1_reg[15]) );
  EDFFX1 \data1_reg_reg[14]  ( .D(data1[14]), .E(n6), .CK(clk), .Q(
        data1_reg[14]) );
  EDFFX1 \data1_reg_reg[13]  ( .D(data1[13]), .E(n7), .CK(clk), .Q(
        data1_reg[13]) );
  EDFFX1 \data1_reg_reg[12]  ( .D(data1[12]), .E(n7), .CK(clk), .Q(
        data1_reg[12]) );
  EDFFX1 \data1_reg_reg[11]  ( .D(data1[11]), .E(n7), .CK(clk), .Q(
        data1_reg[11]) );
  EDFFX1 \data1_reg_reg[10]  ( .D(data1[10]), .E(n7), .CK(clk), .Q(
        data1_reg[10]) );
  EDFFX1 \data1_reg_reg[9]  ( .D(data1[9]), .E(n8), .CK(clk), .Q(data1_reg[9])
         );
  EDFFX1 \data1_reg_reg[8]  ( .D(data1[8]), .E(n8), .CK(clk), .Q(data1_reg[8])
         );
  EDFFX1 \data1_reg_reg[7]  ( .D(data1[7]), .E(n8), .CK(clk), .Q(data1_reg[7])
         );
  EDFFX1 \data1_reg_reg[6]  ( .D(data1[6]), .E(n9), .CK(clk), .Q(data1_reg[6])
         );
  EDFFX1 \data1_reg_reg[5]  ( .D(data1[5]), .E(n14), .CK(clk), .Q(data1_reg[5]) );
  EDFFX1 \data1_reg_reg[4]  ( .D(data1[4]), .E(n14), .CK(clk), .Q(data1_reg[4]) );
  EDFFX1 \data1_reg_reg[3]  ( .D(data1[3]), .E(n13), .CK(clk), .Q(data1_reg[3]) );
  EDFFX1 \data1_reg_reg[2]  ( .D(data1[2]), .E(n9), .CK(clk), .Q(data1_reg[2])
         );
  EDFFX1 \data1_reg_reg[1]  ( .D(data1[1]), .E(n9), .CK(clk), .Q(data1_reg[1])
         );
  EDFFX1 \data1_reg_reg[0]  ( .D(data1[0]), .E(n10), .CK(clk), .Q(data1_reg[0]) );
  EDFFX1 \data2_reg_reg[31]  ( .D(data2[31]), .E(n3), .CK(clk), .Q(
        data2_reg[31]) );
  EDFFX1 \data2_reg_reg[30]  ( .D(data2[30]), .E(n3), .CK(clk), .Q(
        data2_reg[30]) );
  EDFFX1 \data2_reg_reg[29]  ( .D(data2[29]), .E(n3), .CK(clk), .Q(
        data2_reg[29]) );
  EDFFX1 \data2_reg_reg[28]  ( .D(data2[28]), .E(n3), .CK(clk), .Q(
        data2_reg[28]) );
  EDFFX1 \data2_reg_reg[27]  ( .D(data2[27]), .E(n4), .CK(clk), .Q(
        data2_reg[27]) );
  EDFFX1 \data2_reg_reg[26]  ( .D(data2[26]), .E(n4), .CK(clk), .Q(
        data2_reg[26]) );
  EDFFX1 \data2_reg_reg[25]  ( .D(data2[25]), .E(n4), .CK(clk), .Q(
        data2_reg[25]) );
  EDFFX1 \data2_reg_reg[24]  ( .D(data2[24]), .E(n4), .CK(clk), .Q(
        data2_reg[24]) );
  EDFFX1 \data2_reg_reg[23]  ( .D(data2[23]), .E(n4), .CK(clk), .Q(
        data2_reg[23]) );
  EDFFX1 \data2_reg_reg[22]  ( .D(data2[22]), .E(n5), .CK(clk), .Q(
        data2_reg[22]) );
  EDFFX1 \data2_reg_reg[21]  ( .D(data2[21]), .E(n5), .CK(clk), .Q(
        data2_reg[21]) );
  EDFFX1 \data2_reg_reg[20]  ( .D(data2[20]), .E(n5), .CK(clk), .Q(
        data2_reg[20]) );
  EDFFX1 \data2_reg_reg[19]  ( .D(data2[19]), .E(n5), .CK(clk), .Q(
        data2_reg[19]) );
  EDFFX1 \data2_reg_reg[18]  ( .D(data2[18]), .E(n3), .CK(clk), .Q(
        data2_reg[18]) );
  EDFFX1 \data2_reg_reg[17]  ( .D(data2[17]), .E(n6), .CK(clk), .Q(
        data2_reg[17]) );
  EDFFX1 \data2_reg_reg[16]  ( .D(data2[16]), .E(n6), .CK(clk), .Q(
        data2_reg[16]) );
  EDFFX1 \data2_reg_reg[15]  ( .D(data2[15]), .E(n6), .CK(clk), .Q(
        data2_reg[15]) );
  EDFFX1 \data2_reg_reg[14]  ( .D(data2[14]), .E(n6), .CK(clk), .Q(
        data2_reg[14]) );
  EDFFX1 \data2_reg_reg[13]  ( .D(data2[13]), .E(n7), .CK(clk), .Q(
        data2_reg[13]) );
  EDFFX1 \data2_reg_reg[12]  ( .D(data2[12]), .E(n7), .CK(clk), .Q(
        data2_reg[12]) );
  EDFFX1 \data2_reg_reg[11]  ( .D(data2[11]), .E(n7), .CK(clk), .Q(
        data2_reg[11]) );
  EDFFX1 \data2_reg_reg[10]  ( .D(data2[10]), .E(n7), .CK(clk), .Q(
        data2_reg[10]) );
  EDFFX1 \data2_reg_reg[9]  ( .D(data2[9]), .E(n8), .CK(clk), .Q(data2_reg[9])
         );
  EDFFX1 \data2_reg_reg[8]  ( .D(data2[8]), .E(n8), .CK(clk), .Q(data2_reg[8])
         );
  EDFFX1 \data2_reg_reg[7]  ( .D(data2[7]), .E(n8), .CK(clk), .Q(data2_reg[7])
         );
  EDFFX1 \data2_reg_reg[6]  ( .D(data2[6]), .E(n9), .CK(clk), .Q(data2_reg[6])
         );
  EDFFX1 \data2_reg_reg[5]  ( .D(data2[5]), .E(n9), .CK(clk), .Q(data2_reg[5])
         );
  EDFFX1 \data2_reg_reg[4]  ( .D(data2[4]), .E(n9), .CK(clk), .Q(data2_reg[4])
         );
  EDFFX1 \data2_reg_reg[3]  ( .D(data2[3]), .E(n9), .CK(clk), .Q(data2_reg[3])
         );
  EDFFX1 \data2_reg_reg[2]  ( .D(data2[2]), .E(n9), .CK(clk), .Q(data2_reg[2])
         );
  EDFFX1 \data2_reg_reg[1]  ( .D(data2[1]), .E(n14), .CK(clk), .Q(data2_reg[1]) );
  EDFFX1 \data2_reg_reg[0]  ( .D(data2[0]), .E(n14), .CK(clk), .Q(data2_reg[0]) );
  EDFFX1 \sign_extend_reg_reg[31]  ( .D(sign_extend[31]), .E(n11), .CK(clk), 
        .Q(sign_extend_reg[31]) );
  EDFFX1 \sign_extend_reg_reg[30]  ( .D(sign_extend[30]), .E(n11), .CK(clk), 
        .Q(sign_extend_reg[30]) );
  EDFFX1 \sign_extend_reg_reg[29]  ( .D(sign_extend[29]), .E(n11), .CK(clk), 
        .Q(sign_extend_reg[29]) );
  EDFFX1 \sign_extend_reg_reg[28]  ( .D(sign_extend[28]), .E(n11), .CK(clk), 
        .Q(sign_extend_reg[28]) );
  EDFFX1 \sign_extend_reg_reg[27]  ( .D(sign_extend[27]), .E(n11), .CK(clk), 
        .Q(sign_extend_reg[27]) );
  EDFFX1 \sign_extend_reg_reg[26]  ( .D(sign_extend[26]), .E(n11), .CK(clk), 
        .Q(sign_extend_reg[26]) );
  EDFFX1 \sign_extend_reg_reg[25]  ( .D(sign_extend[25]), .E(n12), .CK(clk), 
        .Q(sign_extend_reg[25]) );
  EDFFX1 \sign_extend_reg_reg[24]  ( .D(sign_extend[24]), .E(n12), .CK(clk), 
        .Q(sign_extend_reg[24]) );
  EDFFX1 \sign_extend_reg_reg[23]  ( .D(sign_extend[23]), .E(n12), .CK(clk), 
        .Q(sign_extend_reg[23]) );
  EDFFX1 \sign_extend_reg_reg[22]  ( .D(sign_extend[22]), .E(n12), .CK(clk), 
        .Q(sign_extend_reg[22]) );
  EDFFX1 \sign_extend_reg_reg[21]  ( .D(sign_extend[21]), .E(n12), .CK(clk), 
        .Q(sign_extend_reg[21]) );
  EDFFX1 \sign_extend_reg_reg[20]  ( .D(sign_extend[20]), .E(n12), .CK(clk), 
        .Q(sign_extend_reg[20]) );
  EDFFX1 \sign_extend_reg_reg[19]  ( .D(sign_extend[19]), .E(n12), .CK(clk), 
        .Q(sign_extend_reg[19]) );
  EDFFX1 \sign_extend_reg_reg[18]  ( .D(sign_extend[18]), .E(n12), .CK(clk), 
        .Q(sign_extend_reg[18]) );
  EDFFX1 \sign_extend_reg_reg[17]  ( .D(sign_extend[17]), .E(n12), .CK(clk), 
        .Q(sign_extend_reg[17]) );
  EDFFX1 \sign_extend_reg_reg[16]  ( .D(sign_extend[16]), .E(n12), .CK(clk), 
        .Q(sign_extend_reg[16]) );
  EDFFX1 \sign_extend_reg_reg[15]  ( .D(sign_extend[15]), .E(n12), .CK(clk), 
        .Q(sign_extend_reg[15]) );
  EDFFX1 \sign_extend_reg_reg[14]  ( .D(sign_extend[14]), .E(n12), .CK(clk), 
        .Q(sign_extend_reg[14]) );
  EDFFX1 \sign_extend_reg_reg[13]  ( .D(sign_extend[13]), .E(n13), .CK(clk), 
        .Q(sign_extend_reg[13]) );
  EDFFX1 \sign_extend_reg_reg[12]  ( .D(sign_extend[12]), .E(n13), .CK(clk), 
        .Q(sign_extend_reg[12]) );
  EDFFX1 \sign_extend_reg_reg[11]  ( .D(sign_extend[11]), .E(n13), .CK(clk), 
        .Q(sign_extend_reg[11]) );
  EDFFX1 \sign_extend_reg_reg[10]  ( .D(sign_extend[10]), .E(n13), .CK(clk), 
        .Q(sign_extend_reg[10]) );
  EDFFX1 \sign_extend_reg_reg[9]  ( .D(sign_extend[9]), .E(n7), .CK(clk), .Q(
        sign_extend_reg[9]) );
  EDFFX1 \sign_extend_reg_reg[8]  ( .D(sign_extend[8]), .E(n8), .CK(clk), .Q(
        sign_extend_reg[8]) );
  EDFFX1 \sign_extend_reg_reg[7]  ( .D(sign_extend[7]), .E(n8), .CK(clk), .Q(
        sign_extend_reg[7]) );
  EDFFX1 \sign_extend_reg_reg[6]  ( .D(sign_extend[6]), .E(n8), .CK(clk), .Q(
        sign_extend_reg[6]) );
  EDFFX1 \WB_reg_reg[0]  ( .D(WB[0]), .E(n14), .CK(clk), .Q(WB_reg[0]) );
  EDFFX1 \EX_reg_reg[5]  ( .D(EX[5]), .E(n14), .CK(clk), .Q(EX_reg[5]) );
  EDFFX1 \M_reg_reg[2]  ( .D(M[2]), .E(n10), .CK(clk), .Q(M_reg[2]) );
  EDFFX1 \sign_extend_reg_reg[4]  ( .D(sign_extend[4]), .E(n14), .CK(clk), .Q(
        sign_extend_reg[4]) );
  EDFFX1 \RegRs_reg_reg[0]  ( .D(RegRs[0]), .E(n11), .CK(clk), .Q(RegRs_reg[0]) );
  EDFFX1 \RegRs_reg_reg[2]  ( .D(RegRs[2]), .E(n10), .CK(clk), .Q(RegRs_reg[2]) );
  EDFFX1 \RegRs_reg_reg[1]  ( .D(RegRs[1]), .E(n10), .CK(clk), .Q(RegRs_reg[1]) );
  EDFFX1 \RegRs_reg_reg[4]  ( .D(RegRs[4]), .E(n13), .CK(clk), .Q(RegRs_reg[4]) );
  EDFFX1 \RegRs_reg_reg[3]  ( .D(RegRs[3]), .E(n10), .CK(clk), .Q(RegRs_reg[3]) );
  EDFFX1 \RegRd_reg_reg[4]  ( .D(RegRd[4]), .E(n11), .CK(clk), .Q(RegRd_reg[4]) );
  EDFFX1 \RegRd_reg_reg[2]  ( .D(RegRd[2]), .E(n13), .CK(clk), .Q(RegRd_reg[2]) );
  EDFFX1 \sign_extend_reg_reg[3]  ( .D(sign_extend[3]), .E(n13), .CK(clk), .Q(
        sign_extend_reg[3]) );
  EDFFX1 \RegRd_reg_reg[3]  ( .D(RegRd[3]), .E(n12), .CK(clk), .Q(RegRd_reg[3]) );
  EDFFX1 \RegRd_reg_reg[1]  ( .D(RegRd[1]), .E(n13), .CK(clk), .Q(RegRd_reg[1]) );
  EDFFX1 \RegRd_reg_reg[0]  ( .D(RegRd[0]), .E(n13), .CK(clk), .Q(RegRd_reg[0]) );
  EDFFX1 \sign_extend_reg_reg[2]  ( .D(sign_extend[2]), .E(n13), .CK(clk), .Q(
        sign_extend_reg[2]) );
  EDFFX1 \sign_extend_reg_reg[5]  ( .D(sign_extend[5]), .E(n9), .CK(clk), .Q(
        sign_extend_reg[5]) );
  EDFFX1 \sign_extend_reg_reg[1]  ( .D(sign_extend[1]), .E(n13), .CK(clk), .Q(
        sign_extend_reg[1]) );
  EDFFX1 \RegRt_reg_reg[4]  ( .D(RegRt[4]), .E(n11), .CK(clk), .Q(RegRt_reg[4]) );
  EDFFX1 \RegRt_reg_reg[2]  ( .D(RegRt[2]), .E(n11), .CK(clk), .Q(RegRt_reg[2]) );
  EDFFX1 \RegRt_reg_reg[1]  ( .D(RegRt[1]), .E(n11), .CK(clk), .Q(RegRt_reg[1]) );
  EDFFX1 \RegRt_reg_reg[0]  ( .D(RegRt[0]), .E(n11), .CK(clk), .Q(RegRt_reg[0]) );
  EDFFX1 \RegRt_reg_reg[3]  ( .D(RegRt[3]), .E(n11), .CK(clk), .Q(RegRt_reg[3]) );
  EDFFX1 \sign_extend_reg_reg[0]  ( .D(sign_extend[0]), .E(n13), .CK(clk), .Q(
        sign_extend_reg[0]) );
  EDFFX1 \WB_reg_reg[2]  ( .D(WB[2]), .E(n14), .CK(clk), .Q(WB_reg[2]) );
  EDFFX1 \M_reg_reg[1]  ( .D(M[1]), .E(n14), .CK(clk), .Q(M_reg[1]) );
  EDFFX1 \WB_reg_reg[1]  ( .D(WB[1]), .E(n10), .CK(clk), .Q(WB_reg[1]) );
  EDFFX1 \M_reg_reg[0]  ( .D(M[0]), .E(n10), .CK(clk), .Q(M_reg[0]) );
  EDFFX1 \EX_pcplus4_reg[31]  ( .D(PC_plus4Reg[31]), .E(n3), .CK(clk), .Q(
        EX_pcplus4[31]) );
  EDFFX1 \EX_pcplus4_reg[30]  ( .D(PC_plus4Reg[30]), .E(n3), .CK(clk), .Q(
        EX_pcplus4[30]) );
  EDFFX1 \EX_pcplus4_reg[29]  ( .D(PC_plus4Reg[29]), .E(n3), .CK(clk), .Q(
        EX_pcplus4[29]) );
  EDFFX1 \EX_pcplus4_reg[28]  ( .D(PC_plus4Reg[28]), .E(n3), .CK(clk), .Q(
        EX_pcplus4[28]) );
  EDFFX1 \EX_pcplus4_reg[27]  ( .D(PC_plus4Reg[27]), .E(n4), .CK(clk), .Q(
        EX_pcplus4[27]) );
  EDFFX1 \EX_pcplus4_reg[26]  ( .D(PC_plus4Reg[26]), .E(n4), .CK(clk), .Q(
        EX_pcplus4[26]) );
  EDFFX1 \EX_pcplus4_reg[25]  ( .D(PC_plus4Reg[25]), .E(n4), .CK(clk), .Q(
        EX_pcplus4[25]) );
  EDFFX1 \EX_pcplus4_reg[24]  ( .D(PC_plus4Reg[24]), .E(n4), .CK(clk), .Q(
        EX_pcplus4[24]) );
  EDFFX1 \EX_pcplus4_reg[23]  ( .D(PC_plus4Reg[23]), .E(n5), .CK(clk), .Q(
        EX_pcplus4[23]) );
  EDFFX1 \EX_pcplus4_reg[22]  ( .D(PC_plus4Reg[22]), .E(n5), .CK(clk), .Q(
        EX_pcplus4[22]) );
  EDFFX1 \EX_pcplus4_reg[21]  ( .D(PC_plus4Reg[21]), .E(n5), .CK(clk), .Q(
        EX_pcplus4[21]) );
  EDFFX1 \EX_pcplus4_reg[20]  ( .D(PC_plus4Reg[20]), .E(n5), .CK(clk), .Q(
        EX_pcplus4[20]) );
  EDFFX1 \EX_pcplus4_reg[19]  ( .D(PC_plus4Reg[19]), .E(n6), .CK(clk), .Q(
        EX_pcplus4[19]) );
  EDFFX1 \EX_pcplus4_reg[18]  ( .D(PC_plus4Reg[18]), .E(n6), .CK(clk), .Q(
        EX_pcplus4[18]) );
  EDFFX1 \EX_pcplus4_reg[17]  ( .D(PC_plus4Reg[17]), .E(n6), .CK(clk), .Q(
        EX_pcplus4[17]) );
  EDFFX1 \EX_pcplus4_reg[16]  ( .D(PC_plus4Reg[16]), .E(n6), .CK(clk), .Q(
        EX_pcplus4[16]) );
  EDFFX1 \EX_pcplus4_reg[15]  ( .D(PC_plus4Reg[15]), .E(n6), .CK(clk), .Q(
        EX_pcplus4[15]) );
  EDFFX1 \EX_pcplus4_reg[14]  ( .D(PC_plus4Reg[14]), .E(n7), .CK(clk), .Q(
        EX_pcplus4[14]) );
  EDFFX1 \EX_pcplus4_reg[13]  ( .D(PC_plus4Reg[13]), .E(n7), .CK(clk), .Q(
        EX_pcplus4[13]) );
  EDFFX1 \EX_pcplus4_reg[12]  ( .D(PC_plus4Reg[12]), .E(n7), .CK(clk), .Q(
        EX_pcplus4[12]) );
  EDFFX1 \EX_pcplus4_reg[11]  ( .D(PC_plus4Reg[11]), .E(n7), .CK(clk), .Q(
        EX_pcplus4[11]) );
  EDFFX1 \EX_pcplus4_reg[10]  ( .D(PC_plus4Reg[10]), .E(n8), .CK(clk), .Q(
        EX_pcplus4[10]) );
  EDFFX1 \EX_pcplus4_reg[9]  ( .D(PC_plus4Reg[9]), .E(n8), .CK(clk), .Q(
        EX_pcplus4[9]) );
  EDFFX1 \EX_pcplus4_reg[8]  ( .D(PC_plus4Reg[8]), .E(n8), .CK(clk), .Q(
        EX_pcplus4[8]) );
  EDFFX1 \EX_pcplus4_reg[7]  ( .D(PC_plus4Reg[7]), .E(n8), .CK(clk), .Q(
        EX_pcplus4[7]) );
  EDFFX1 \EX_pcplus4_reg[6]  ( .D(PC_plus4Reg[6]), .E(n10), .CK(clk), .Q(
        EX_pcplus4[6]) );
  EDFFX1 \EX_pcplus4_reg[5]  ( .D(PC_plus4Reg[5]), .E(n10), .CK(clk), .Q(
        EX_pcplus4[5]) );
  EDFFX1 \EX_pcplus4_reg[4]  ( .D(PC_plus4Reg[4]), .E(n10), .CK(clk), .Q(
        EX_pcplus4[4]) );
  EDFFX1 \EX_pcplus4_reg[3]  ( .D(PC_plus4Reg[3]), .E(n10), .CK(clk), .Q(
        EX_pcplus4[3]) );
  EDFFX1 \EX_pcplus4_reg[2]  ( .D(PC_plus4Reg[2]), .E(n10), .CK(clk), .Q(
        EX_pcplus4[2]) );
  EDFFX1 \EX_pcplus4_reg[1]  ( .D(PC_plus4Reg[1]), .E(n14), .CK(clk), .Q(
        EX_pcplus4[1]) );
  EDFFX1 \EX_pcplus4_reg[0]  ( .D(PC_plus4Reg[0]), .E(n14), .CK(clk), .Q(
        EX_pcplus4[0]) );
  EDFFX1 \EX_reg_reg[3]  ( .D(EX[3]), .E(n9), .CK(clk), .QN(n1) );
  INVX6 U2 ( .A(n1), .Y(EX_reg[3]) );
  CLKBUFX3 U3 ( .A(n4), .Y(n10) );
  CLKBUFX3 U4 ( .A(n8), .Y(n6) );
  CLKBUFX3 U5 ( .A(n8), .Y(n5) );
  CLKBUFX3 U6 ( .A(stall_bothzero), .Y(n4) );
  CLKBUFX3 U7 ( .A(n4), .Y(n3) );
  CLKBUFX3 U8 ( .A(n4), .Y(n9) );
  CLKBUFX3 U9 ( .A(stall_bothzero), .Y(n8) );
  CLKBUFX3 U10 ( .A(n8), .Y(n7) );
  CLKBUFX3 U11 ( .A(n4), .Y(n13) );
  CLKBUFX3 U12 ( .A(n4), .Y(n12) );
  CLKBUFX3 U13 ( .A(n8), .Y(n11) );
  CLKBUFX3 U14 ( .A(n8), .Y(n14) );
endmodule


module ALUcontrol ( ALUctrl, ALUOp, func_field );
  output [3:0] ALUctrl;
  input [2:0] ALUOp;
  input [5:0] func_field;
  wire   n19, n20, n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;

  CLKMX2X2 U1 ( .A(n5), .B(n6), .S0(func_field[0]), .Y(n1) );
  INVX6 U2 ( .A(n1), .Y(ALUctrl[3]) );
  NAND2X6 U3 ( .A(n7), .B(n8), .Y(ALUctrl[2]) );
  MX2XL U4 ( .A(n6), .B(n5), .S0(func_field[0]), .Y(n7) );
  CLKBUFX6 U5 ( .A(n19), .Y(ALUctrl[1]) );
  BUFX12 U6 ( .A(n20), .Y(ALUctrl[0]) );
  NAND4BXL U7 ( .AN(n16), .B(func_field[5]), .C(func_field[1]), .D(n17), .Y(n8) );
  NOR2BX1 U8 ( .AN(n6), .B(n9), .Y(n19) );
  NAND2X1 U9 ( .A(func_field[1]), .B(n10), .Y(n6) );
  OAI21XL U10 ( .A0(n8), .A1(n11), .B0(n12), .Y(n20) );
  MXI2X1 U11 ( .A(n13), .B(n9), .S0(func_field[0]), .Y(n12) );
  OAI21XL U12 ( .A0(func_field[1]), .A1(n14), .B0(n5), .Y(n13) );
  NAND2X1 U13 ( .A(n9), .B(func_field[1]), .Y(n5) );
  AND3X1 U14 ( .A(func_field[2]), .B(n15), .C(func_field[5]), .Y(n9) );
  CLKINVX1 U15 ( .A(n10), .Y(n14) );
  NOR3BXL U16 ( .AN(n15), .B(func_field[2]), .C(func_field[5]), .Y(n10) );
  NOR2X1 U17 ( .A(n16), .B(func_field[3]), .Y(n15) );
  CLKINVX1 U18 ( .A(func_field[3]), .Y(n11) );
  NOR2X1 U19 ( .A(func_field[2]), .B(func_field[0]), .Y(n17) );
  NAND3BX1 U20 ( .AN(ALUOp[0]), .B(ALUOp[1]), .C(n18), .Y(n16) );
  NOR2X1 U21 ( .A(func_field[4]), .B(ALUOp[2]), .Y(n18) );
endmodule


module fowarding_unit ( ID_EX_Rs, ID_EX_Rt, EX_MEM_RegWrite, MEM_WB_RegWrite, 
        EX_MEM_Rd, MEM_WB_Rd, Foward_A, Foward_B );
  input [4:0] ID_EX_Rs;
  input [4:0] ID_EX_Rt;
  input [4:0] EX_MEM_Rd;
  input [4:0] MEM_WB_Rd;
  output [1:0] Foward_A;
  output [1:0] Foward_B;
  input EX_MEM_RegWrite, MEM_WB_RegWrite;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;

  NOR2X1 U1 ( .A(Foward_A[1]), .B(n1), .Y(Foward_B[1]) );
  NOR4X1 U2 ( .A(n2), .B(n3), .C(n4), .D(n5), .Y(Foward_B[0]) );
  XOR2X1 U3 ( .A(MEM_WB_Rd[2]), .B(ID_EX_Rt[2]), .Y(n5) );
  XOR2X1 U4 ( .A(MEM_WB_Rd[1]), .B(ID_EX_Rt[1]), .Y(n4) );
  XOR2X1 U5 ( .A(MEM_WB_Rd[4]), .B(ID_EX_Rt[4]), .Y(n3) );
  NAND4BX1 U6 ( .AN(n6), .B(n7), .C(n8), .D(n9), .Y(n2) );
  XNOR2X1 U7 ( .A(ID_EX_Rt[3]), .B(MEM_WB_Rd[3]), .Y(n8) );
  XNOR2X1 U8 ( .A(ID_EX_Rt[0]), .B(MEM_WB_Rd[0]), .Y(n7) );
  CLKINVX1 U9 ( .A(n10), .Y(Foward_A[1]) );
  NOR2X1 U10 ( .A(n6), .B(n9), .Y(Foward_A[0]) );
  NAND4X1 U11 ( .A(n11), .B(n12), .C(n13), .D(n14), .Y(n9) );
  XNOR2X1 U12 ( .A(ID_EX_Rs[1]), .B(MEM_WB_Rd[1]), .Y(n14) );
  NOR2X1 U13 ( .A(n15), .B(n16), .Y(n13) );
  XOR2X1 U14 ( .A(MEM_WB_Rd[0]), .B(ID_EX_Rs[0]), .Y(n16) );
  XOR2X1 U15 ( .A(MEM_WB_Rd[2]), .B(ID_EX_Rs[2]), .Y(n15) );
  XNOR2X1 U16 ( .A(ID_EX_Rs[3]), .B(MEM_WB_Rd[3]), .Y(n12) );
  XNOR2X1 U17 ( .A(ID_EX_Rs[4]), .B(MEM_WB_Rd[4]), .Y(n11) );
  NAND4X1 U18 ( .A(MEM_WB_RegWrite), .B(n17), .C(n1), .D(n10), .Y(n6) );
  NAND4X1 U19 ( .A(n18), .B(n19), .C(n20), .D(n21), .Y(n10) );
  NOR3X1 U20 ( .A(n22), .B(n23), .C(n24), .Y(n21) );
  XOR2X1 U21 ( .A(ID_EX_Rs[2]), .B(EX_MEM_Rd[2]), .Y(n24) );
  XOR2X1 U22 ( .A(ID_EX_Rs[4]), .B(EX_MEM_Rd[4]), .Y(n23) );
  XOR2X1 U23 ( .A(ID_EX_Rs[3]), .B(EX_MEM_Rd[3]), .Y(n22) );
  XNOR2X1 U24 ( .A(EX_MEM_Rd[0]), .B(ID_EX_Rs[0]), .Y(n20) );
  XNOR2X1 U25 ( .A(EX_MEM_Rd[1]), .B(ID_EX_Rs[1]), .Y(n18) );
  NAND4X1 U26 ( .A(n25), .B(n19), .C(n26), .D(n27), .Y(n1) );
  NOR3X1 U27 ( .A(n28), .B(n29), .C(n30), .Y(n27) );
  XOR2X1 U28 ( .A(ID_EX_Rt[2]), .B(EX_MEM_Rd[2]), .Y(n30) );
  XOR2X1 U29 ( .A(ID_EX_Rt[4]), .B(EX_MEM_Rd[4]), .Y(n29) );
  XOR2X1 U30 ( .A(ID_EX_Rt[3]), .B(EX_MEM_Rd[3]), .Y(n28) );
  XNOR2X1 U31 ( .A(EX_MEM_Rd[0]), .B(ID_EX_Rt[0]), .Y(n26) );
  CLKINVX1 U32 ( .A(n31), .Y(n19) );
  OAI31XL U33 ( .A0(n32), .A1(EX_MEM_Rd[1]), .A2(EX_MEM_Rd[0]), .B0(
        EX_MEM_RegWrite), .Y(n31) );
  OR3X1 U34 ( .A(EX_MEM_Rd[3]), .B(EX_MEM_Rd[4]), .C(EX_MEM_Rd[2]), .Y(n32) );
  XNOR2X1 U35 ( .A(EX_MEM_Rd[1]), .B(ID_EX_Rt[1]), .Y(n25) );
  OR4X1 U36 ( .A(MEM_WB_Rd[0]), .B(MEM_WB_Rd[1]), .C(n33), .D(MEM_WB_Rd[2]), 
        .Y(n17) );
  OR2X1 U37 ( .A(MEM_WB_Rd[4]), .B(MEM_WB_Rd[3]), .Y(n33) );
endmodule


module alu_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [32:0] carry;
  wire   [31:0] B_AS;
  assign carry[0] = ADD_SUB;

  ADDFXL U1_30 ( .A(A[30]), .B(B_AS[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B_AS[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B_AS[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B_AS[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B_AS[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B_AS[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B_AS[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B_AS[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B_AS[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B_AS[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B_AS[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B_AS[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B_AS[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B_AS[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B_AS[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B_AS[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B_AS[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B_AS[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B_AS[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B_AS[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B_AS[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B_AS[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B_AS[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B_AS[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B_AS[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B_AS[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B_AS[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDFXL U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(carry[0]), .CO(carry[1]), .S(SUM[0]) );
  XOR3XL U1_31 ( .A(A[31]), .B(B_AS[31]), .C(carry[31]), .Y(SUM[31]) );
  XOR2X1 U1 ( .A(B[9]), .B(carry[0]), .Y(B_AS[9]) );
  XOR2X1 U2 ( .A(B[8]), .B(carry[0]), .Y(B_AS[8]) );
  XOR2X1 U3 ( .A(B[7]), .B(carry[0]), .Y(B_AS[7]) );
  XOR2X1 U4 ( .A(B[6]), .B(carry[0]), .Y(B_AS[6]) );
  XOR2X1 U5 ( .A(B[5]), .B(carry[0]), .Y(B_AS[5]) );
  XOR2X1 U6 ( .A(B[4]), .B(carry[0]), .Y(B_AS[4]) );
  XOR2X1 U7 ( .A(B[3]), .B(carry[0]), .Y(B_AS[3]) );
  XOR2X1 U8 ( .A(B[31]), .B(carry[0]), .Y(B_AS[31]) );
  XOR2X1 U9 ( .A(B[30]), .B(carry[0]), .Y(B_AS[30]) );
  XOR2X1 U10 ( .A(B[2]), .B(carry[0]), .Y(B_AS[2]) );
  XOR2X1 U11 ( .A(B[29]), .B(carry[0]), .Y(B_AS[29]) );
  XOR2X1 U12 ( .A(B[28]), .B(carry[0]), .Y(B_AS[28]) );
  XOR2X1 U13 ( .A(B[27]), .B(carry[0]), .Y(B_AS[27]) );
  XOR2X1 U14 ( .A(B[26]), .B(carry[0]), .Y(B_AS[26]) );
  XOR2X1 U15 ( .A(B[25]), .B(carry[0]), .Y(B_AS[25]) );
  XOR2X1 U16 ( .A(B[24]), .B(carry[0]), .Y(B_AS[24]) );
  XOR2X1 U17 ( .A(B[23]), .B(carry[0]), .Y(B_AS[23]) );
  XOR2X1 U18 ( .A(B[22]), .B(carry[0]), .Y(B_AS[22]) );
  XOR2X1 U19 ( .A(B[21]), .B(carry[0]), .Y(B_AS[21]) );
  XOR2X1 U20 ( .A(B[20]), .B(carry[0]), .Y(B_AS[20]) );
  XOR2X1 U21 ( .A(B[1]), .B(carry[0]), .Y(B_AS[1]) );
  XOR2X1 U22 ( .A(B[19]), .B(carry[0]), .Y(B_AS[19]) );
  XOR2X1 U23 ( .A(B[18]), .B(carry[0]), .Y(B_AS[18]) );
  XOR2X1 U24 ( .A(B[17]), .B(carry[0]), .Y(B_AS[17]) );
  XOR2X1 U25 ( .A(B[16]), .B(carry[0]), .Y(B_AS[16]) );
  XOR2X1 U26 ( .A(B[15]), .B(carry[0]), .Y(B_AS[15]) );
  XOR2X1 U27 ( .A(B[14]), .B(carry[0]), .Y(B_AS[14]) );
  XOR2X1 U28 ( .A(B[13]), .B(carry[0]), .Y(B_AS[13]) );
  XOR2X1 U29 ( .A(B[12]), .B(carry[0]), .Y(B_AS[12]) );
  XOR2X1 U30 ( .A(B[11]), .B(carry[0]), .Y(B_AS[11]) );
  XOR2X1 U31 ( .A(B[10]), .B(carry[0]), .Y(B_AS[10]) );
  XOR2X1 U32 ( .A(B[0]), .B(carry[0]), .Y(B_AS[0]) );
endmodule


module alu_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104;

  INVXL U1 ( .A(B[2]), .Y(n15) );
  INVXL U2 ( .A(B[3]), .Y(n17) );
  INVXL U3 ( .A(B[27]), .Y(n12) );
  INVXL U4 ( .A(B[20]), .Y(n8) );
  INVXL U5 ( .A(B[21]), .Y(n9) );
  INVXL U6 ( .A(B[28]), .Y(n13) );
  INVX1 U7 ( .A(B[29]), .Y(n14) );
  INVXL U8 ( .A(B[26]), .Y(n11) );
  INVXL U9 ( .A(B[9]), .Y(n20) );
  INVXL U10 ( .A(B[19]), .Y(n6) );
  NOR2XL U11 ( .A(n29), .B(B[4]), .Y(n104) );
  NOR2BXL U12 ( .AN(A[5]), .B(B[5]), .Y(n98) );
  NAND2XL U13 ( .A(A[9]), .B(n20), .Y(n91) );
  NAND2XL U14 ( .A(A[12]), .B(n3), .Y(n84) );
  NAND2XL U15 ( .A(A[21]), .B(n9), .Y(n53) );
  NAND2XL U16 ( .A(A[13]), .B(n4), .Y(n81) );
  NAND2XL U17 ( .A(A[20]), .B(n8), .Y(n52) );
  NAND2XL U18 ( .A(A[10]), .B(n1), .Y(n90) );
  NAND2XL U19 ( .A(A[11]), .B(n2), .Y(n85) );
  NAND2XL U20 ( .A(A[29]), .B(n14), .Y(n37) );
  NAND2XL U21 ( .A(A[28]), .B(n13), .Y(n39) );
  NAND2XL U22 ( .A(A[27]), .B(n12), .Y(n43) );
  NAND2XL U23 ( .A(A[26]), .B(n11), .Y(n44) );
  NAND2XL U24 ( .A(A[19]), .B(n6), .Y(n47) );
  NAND2XL U25 ( .A(A[3]), .B(n17), .Y(n60) );
  NAND2XL U26 ( .A(A[2]), .B(n15), .Y(n59) );
  NAND2BXL U27 ( .AN(A[5]), .B(B[5]), .Y(n97) );
  NOR2XL U28 ( .A(A[19]), .B(n6), .Y(n73) );
  OAI32XL U29 ( .A0(n75), .A1(n49), .A2(n50), .B0(A[18]), .B1(n5), .Y(n74) );
  NOR2BXL U30 ( .AN(B[0]), .B(A[0]), .Y(n102) );
  NAND2BXL U31 ( .AN(B[22]), .B(A[22]), .Y(n54) );
  NAND2BXL U32 ( .AN(B[14]), .B(A[14]), .Y(n80) );
  NAND2BXL U33 ( .AN(A[23]), .B(B[23]), .Y(n70) );
  NAND2BXL U34 ( .AN(A[15]), .B(B[15]), .Y(n78) );
  NOR2XL U35 ( .A(A[9]), .B(n20), .Y(n88) );
  NOR2BXL U36 ( .AN(A[18]), .B(B[18]), .Y(n50) );
  NOR2BXL U37 ( .AN(A[31]), .B(B[31]), .Y(n61) );
  NOR2BXL U38 ( .AN(A[15]), .B(B[15]), .Y(n79) );
  NOR2BXL U39 ( .AN(A[23]), .B(B[23]), .Y(n51) );
  NOR2BXL U40 ( .AN(A[8]), .B(B[8]), .Y(n94) );
  OAI32XL U41 ( .A0(n67), .A1(n41), .A2(n10), .B0(A[26]), .B1(n11), .Y(n66) );
  INVXL U42 ( .A(B[1]), .Y(n7) );
  NOR2BXL U43 ( .AN(A[0]), .B(B[0]), .Y(n40) );
  INVXL U44 ( .A(B[11]), .Y(n2) );
  INVXL U45 ( .A(B[13]), .Y(n4) );
  INVXL U46 ( .A(B[10]), .Y(n1) );
  INVXL U47 ( .A(B[12]), .Y(n3) );
  AO21XL U48 ( .A0(n24), .A1(n102), .B0(B[1]), .Y(n103) );
  CLKINVX1 U49 ( .A(n104), .Y(n18) );
  CLKINVX1 U50 ( .A(B[31]), .Y(n16) );
  CLKINVX1 U51 ( .A(B[8]), .Y(n19) );
  INVXL U52 ( .A(A[1]), .Y(n24) );
  INVXL U53 ( .A(A[4]), .Y(n29) );
  INVXL U54 ( .A(A[25]), .Y(n27) );
  INVXL U55 ( .A(A[7]), .Y(n31) );
  INVXL U56 ( .A(A[24]), .Y(n26) );
  INVXL U57 ( .A(A[6]), .Y(n30) );
  INVXL U58 ( .A(A[17]), .Y(n23) );
  INVXL U59 ( .A(A[30]), .Y(n28) );
  INVXL U60 ( .A(A[16]), .Y(n22) );
  INVXL U61 ( .A(A[22]), .Y(n25) );
  INVXL U62 ( .A(A[14]), .Y(n21) );
  CLKINVX1 U63 ( .A(n44), .Y(n10) );
  CLKINVX1 U64 ( .A(B[18]), .Y(n5) );
  NOR4X1 U65 ( .A(n32), .B(n33), .C(n34), .D(n35), .Y(EQ) );
  NAND4X1 U66 ( .A(n36), .B(n37), .C(n38), .D(n39), .Y(n35) );
  OAI22XL U67 ( .A0(A[1]), .A1(n40), .B0(n40), .B1(n7), .Y(n36) );
  NAND4BBXL U68 ( .AN(n41), .BN(n42), .C(n43), .D(n44), .Y(n34) );
  NAND2BX1 U69 ( .AN(n45), .B(n46), .Y(n33) );
  NOR4BX1 U70 ( .AN(n47), .B(n48), .C(n49), .D(n50), .Y(n46) );
  NAND4BX1 U71 ( .AN(n51), .B(n52), .C(n53), .D(n54), .Y(n45) );
  NAND4BBXL U72 ( .AN(n55), .BN(n56), .C(n57), .D(n58), .Y(n32) );
  NOR4BBX1 U73 ( .AN(n59), .BN(n60), .C(LT), .D(n61), .Y(n58) );
  OAI22XL U74 ( .A0(A[31]), .A1(n16), .B0(n61), .B1(n62), .Y(LT) );
  AOI32X1 U75 ( .A0(n37), .A1(n38), .A2(n63), .B0(B[30]), .B1(n28), .Y(n62) );
  OAI221XL U76 ( .A0(A[28]), .A1(n13), .B0(A[29]), .B1(n14), .C0(n64), .Y(n63)
         );
  OAI211X1 U77 ( .A0(n65), .A1(n66), .B0(n39), .C0(n43), .Y(n64) );
  NOR2X1 U78 ( .A(n27), .B(B[25]), .Y(n41) );
  AOI221XL U79 ( .A0(B[25]), .A1(n27), .B0(B[24]), .B1(n26), .C0(n68), .Y(n67)
         );
  AOI211X1 U80 ( .A0(n69), .A1(n70), .B0(n51), .C0(n42), .Y(n68) );
  NOR2X1 U81 ( .A(n26), .B(B[24]), .Y(n42) );
  AOI32X1 U82 ( .A0(n54), .A1(n53), .A2(n71), .B0(B[22]), .B1(n25), .Y(n69) );
  OAI221XL U83 ( .A0(A[20]), .A1(n8), .B0(A[21]), .B1(n9), .C0(n72), .Y(n71)
         );
  OAI211X1 U84 ( .A0(n73), .A1(n74), .B0(n52), .C0(n47), .Y(n72) );
  NOR2X1 U85 ( .A(n23), .B(B[17]), .Y(n49) );
  AOI221XL U86 ( .A0(B[17]), .A1(n23), .B0(B[16]), .B1(n22), .C0(n76), .Y(n75)
         );
  AOI211X1 U87 ( .A0(n77), .A1(n78), .B0(n79), .C0(n48), .Y(n76) );
  NOR2X1 U88 ( .A(n22), .B(B[16]), .Y(n48) );
  AOI32X1 U89 ( .A0(n80), .A1(n81), .A2(n82), .B0(B[14]), .B1(n21), .Y(n77) );
  OAI221XL U90 ( .A0(A[12]), .A1(n3), .B0(A[13]), .B1(n4), .C0(n83), .Y(n82)
         );
  NAND3X1 U91 ( .A(n84), .B(n85), .C(n86), .Y(n83) );
  OAI221XL U92 ( .A0(A[10]), .A1(n1), .B0(A[11]), .B1(n2), .C0(n87), .Y(n86)
         );
  OAI211X1 U93 ( .A0(n88), .A1(n89), .B0(n90), .C0(n91), .Y(n87) );
  OAI32X1 U94 ( .A0(n92), .A1(n93), .A2(n94), .B0(A[8]), .B1(n19), .Y(n89) );
  AOI221XL U95 ( .A0(B[7]), .A1(n31), .B0(B[6]), .B1(n30), .C0(n95), .Y(n92)
         );
  AOI211X1 U96 ( .A0(n96), .A1(n97), .B0(n98), .C0(n99), .Y(n95) );
  AOI32X1 U97 ( .A0(n18), .A1(n60), .A2(n100), .B0(B[4]), .B1(n29), .Y(n96) );
  OAI221XL U98 ( .A0(A[2]), .A1(n15), .B0(A[3]), .B1(n17), .C0(n101), .Y(n100)
         );
  OAI211X1 U99 ( .A0(n102), .A1(n24), .B0(n103), .C0(n59), .Y(n101) );
  NOR2X1 U100 ( .A(A[27]), .B(n12), .Y(n65) );
  OR2X1 U101 ( .A(B[30]), .B(n28), .Y(n38) );
  NOR4X1 U102 ( .A(n104), .B(n98), .C(n99), .D(n93), .Y(n57) );
  NOR2X1 U103 ( .A(n31), .B(B[7]), .Y(n93) );
  NOR2X1 U104 ( .A(n30), .B(B[6]), .Y(n99) );
  NAND4BX1 U105 ( .AN(n94), .B(n91), .C(n90), .D(n85), .Y(n56) );
  NAND4BX1 U106 ( .AN(n79), .B(n84), .C(n81), .D(n80), .Y(n55) );
endmodule


module alu_DW_leftsh_1 ( A, SH, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n213, n214, n215,
         n216, n217, n220, n321, n322, n323, n324, n325, n326;

  MXI2XL U255 ( .A(A[17]), .B(A[16]), .S0(SH[0]), .Y(n181) );
  MXI2XL U256 ( .A(A[7]), .B(A[6]), .S0(SH[0]), .Y(n171) );
  MXI2XL U257 ( .A(A[25]), .B(A[24]), .S0(SH[0]), .Y(n189) );
  MXI2XL U258 ( .A(A[18]), .B(A[17]), .S0(SH[0]), .Y(n182) );
  MXI2XL U259 ( .A(A[2]), .B(A[1]), .S0(SH[0]), .Y(n166) );
  MXI2XL U260 ( .A(A[1]), .B(A[0]), .S0(SH[0]), .Y(n165) );
  MXI2XL U261 ( .A(A[12]), .B(A[11]), .S0(SH[0]), .Y(n176) );
  MXI2XL U262 ( .A(A[26]), .B(A[25]), .S0(SH[0]), .Y(n190) );
  MXI2XL U263 ( .A(A[16]), .B(A[15]), .S0(SH[0]), .Y(n180) );
  MXI2XL U264 ( .A(A[15]), .B(A[14]), .S0(SH[0]), .Y(n179) );
  MXI2XL U265 ( .A(A[29]), .B(A[28]), .S0(SH[0]), .Y(n193) );
  MXI2XL U266 ( .A(A[6]), .B(A[5]), .S0(SH[0]), .Y(n170) );
  MXI2XL U267 ( .A(A[5]), .B(A[4]), .S0(SH[0]), .Y(n169) );
  MXI2XL U268 ( .A(A[24]), .B(A[23]), .S0(SH[0]), .Y(n188) );
  MXI2XL U269 ( .A(A[23]), .B(A[22]), .S0(SH[0]), .Y(n187) );
  MXI2XL U270 ( .A(A[20]), .B(A[19]), .S0(SH[0]), .Y(n184) );
  MXI2XL U271 ( .A(A[19]), .B(A[18]), .S0(SH[0]), .Y(n183) );
  MXI2XL U272 ( .A(A[22]), .B(A[21]), .S0(SH[0]), .Y(n186) );
  MXI2XL U273 ( .A(A[21]), .B(A[20]), .S0(SH[0]), .Y(n185) );
  MXI2XL U274 ( .A(A[14]), .B(A[13]), .S0(SH[0]), .Y(n178) );
  MXI2XL U275 ( .A(A[13]), .B(A[12]), .S0(SH[0]), .Y(n177) );
  MXI2XL U276 ( .A(A[11]), .B(A[10]), .S0(SH[0]), .Y(n175) );
  MXI2XL U277 ( .A(A[10]), .B(A[9]), .S0(SH[0]), .Y(n174) );
  MXI2XL U278 ( .A(A[4]), .B(A[3]), .S0(SH[0]), .Y(n168) );
  MXI2XL U279 ( .A(A[3]), .B(A[2]), .S0(SH[0]), .Y(n167) );
  MXI2XL U280 ( .A(A[9]), .B(A[8]), .S0(SH[0]), .Y(n173) );
  MXI2XL U281 ( .A(A[8]), .B(A[7]), .S0(SH[0]), .Y(n172) );
  MXI2XL U282 ( .A(A[28]), .B(A[27]), .S0(SH[0]), .Y(n192) );
  MXI2XL U283 ( .A(A[27]), .B(A[26]), .S0(SH[0]), .Y(n191) );
  MXI2XL U284 ( .A(n116), .B(n108), .S0(SH[3]), .Y(n84) );
  MXI2XL U285 ( .A(n117), .B(n109), .S0(SH[3]), .Y(n85) );
  MXI2XL U286 ( .A(n118), .B(n110), .S0(SH[3]), .Y(n86) );
  MXI2XL U287 ( .A(n119), .B(n111), .S0(SH[3]), .Y(n87) );
  MXI2XL U288 ( .A(n120), .B(n112), .S0(SH[3]), .Y(n88) );
  MXI2XL U289 ( .A(n121), .B(n113), .S0(SH[3]), .Y(n89) );
  MXI2XL U290 ( .A(n122), .B(n114), .S0(SH[3]), .Y(n90) );
  MXI2XL U291 ( .A(n123), .B(n115), .S0(SH[3]), .Y(n91) );
  NOR2XL U292 ( .A(n164), .B(SH[1]), .Y(n132) );
  NOR2XL U293 ( .A(n165), .B(SH[1]), .Y(n133) );
  MXI2XL U294 ( .A(n195), .B(n193), .S0(SH[1]), .Y(n163) );
  NOR2XL U295 ( .A(n102), .B(SH[3]), .Y(n70) );
  NOR2XL U296 ( .A(n103), .B(SH[3]), .Y(n71) );
  NOR2XL U297 ( .A(n104), .B(SH[3]), .Y(n72) );
  NOR2XL U298 ( .A(n105), .B(SH[3]), .Y(n73) );
  NOR2XL U299 ( .A(n106), .B(SH[3]), .Y(n74) );
  NOR2XL U300 ( .A(n107), .B(SH[3]), .Y(n75) );
  NOR2XL U301 ( .A(n101), .B(SH[3]), .Y(n69) );
  NOR2XL U302 ( .A(n100), .B(SH[3]), .Y(n68) );
  MXI2XL U303 ( .A(n128), .B(n120), .S0(SH[3]), .Y(n96) );
  MXI2XL U304 ( .A(n160), .B(n156), .S0(SH[2]), .Y(n128) );
  MXI2XL U305 ( .A(n192), .B(n190), .S0(SH[1]), .Y(n160) );
  MXI2XL U306 ( .A(n129), .B(n121), .S0(SH[3]), .Y(n97) );
  MXI2XL U307 ( .A(n161), .B(n157), .S0(SH[2]), .Y(n129) );
  MXI2XL U308 ( .A(n193), .B(n191), .S0(SH[1]), .Y(n161) );
  MXI2XL U309 ( .A(n130), .B(n122), .S0(SH[3]), .Y(n98) );
  MXI2XL U310 ( .A(n162), .B(n158), .S0(SH[2]), .Y(n130) );
  MXI2XL U311 ( .A(n194), .B(n192), .S0(SH[1]), .Y(n162) );
  MXI2XL U312 ( .A(n124), .B(n116), .S0(SH[3]), .Y(n92) );
  MXI2XL U313 ( .A(n156), .B(n152), .S0(SH[2]), .Y(n124) );
  MXI2XL U314 ( .A(n125), .B(n117), .S0(SH[3]), .Y(n93) );
  MXI2XL U315 ( .A(n157), .B(n153), .S0(SH[2]), .Y(n125) );
  MXI2XL U316 ( .A(n126), .B(n118), .S0(SH[3]), .Y(n94) );
  MXI2XL U317 ( .A(n158), .B(n154), .S0(SH[2]), .Y(n126) );
  MXI2XL U318 ( .A(n127), .B(n119), .S0(SH[3]), .Y(n95) );
  MXI2XL U319 ( .A(n159), .B(n155), .S0(SH[2]), .Y(n127) );
  NOR2XL U320 ( .A(n67), .B(SH[5]), .Y(n35) );
  MXI2XL U321 ( .A(n99), .B(n83), .S0(SH[4]), .Y(n67) );
  MXI2XL U322 ( .A(n131), .B(n123), .S0(SH[3]), .Y(n99) );
  MXI2XL U323 ( .A(n163), .B(n159), .S0(SH[2]), .Y(n131) );
  NOR2XL U324 ( .A(SH[9]), .B(SH[8]), .Y(n321) );
  NOR2XL U325 ( .A(SH[11]), .B(SH[10]), .Y(n322) );
  NOR2XL U326 ( .A(SH[25]), .B(SH[26]), .Y(n323) );
  NOR2XL U327 ( .A(SH[27]), .B(SH[28]), .Y(n324) );
  NOR2XL U328 ( .A(SH[13]), .B(SH[14]), .Y(n325) );
  OR2XL U329 ( .A(SH[19]), .B(SH[20]), .Y(n215) );
  OR2XL U330 ( .A(SH[21]), .B(SH[22]), .Y(n216) );
  OR2XL U331 ( .A(SH[31]), .B(SH[12]), .Y(n208) );
  OR2XL U332 ( .A(SH[29]), .B(SH[30]), .Y(n220) );
  OR2X6 U333 ( .A(n197), .B(n198), .Y(n3) );
  OR2X1 U334 ( .A(n199), .B(n200), .Y(n197) );
  OR2X1 U335 ( .A(n201), .B(n202), .Y(n198) );
  OR2X1 U336 ( .A(n206), .B(n207), .Y(n199) );
  NOR2BX1 U337 ( .AN(n4), .B(n3), .Y(B[0]) );
  NOR2XL U338 ( .A(n36), .B(SH[5]), .Y(n4) );
  NOR2BX1 U339 ( .AN(n6), .B(n3), .Y(B[2]) );
  NOR2XL U340 ( .A(n38), .B(SH[5]), .Y(n6) );
  NAND2BXL U341 ( .AN(SH[4]), .B(n70), .Y(n38) );
  NOR2BX1 U342 ( .AN(n7), .B(n3), .Y(B[3]) );
  NOR2XL U343 ( .A(n39), .B(SH[5]), .Y(n7) );
  NAND2BXL U344 ( .AN(SH[4]), .B(n71), .Y(n39) );
  NOR2BX1 U345 ( .AN(n8), .B(n3), .Y(B[4]) );
  NOR2XL U346 ( .A(n40), .B(SH[5]), .Y(n8) );
  NAND2BXL U347 ( .AN(SH[4]), .B(n72), .Y(n40) );
  NOR2BX1 U348 ( .AN(n9), .B(n3), .Y(B[5]) );
  NOR2XL U349 ( .A(n41), .B(SH[5]), .Y(n9) );
  NAND2BXL U350 ( .AN(SH[4]), .B(n73), .Y(n41) );
  NOR2BX1 U351 ( .AN(n10), .B(n3), .Y(B[6]) );
  NOR2XL U352 ( .A(n42), .B(SH[5]), .Y(n10) );
  NAND2BXL U353 ( .AN(SH[4]), .B(n74), .Y(n42) );
  NOR2BX1 U354 ( .AN(n11), .B(n3), .Y(B[7]) );
  NOR2XL U355 ( .A(n43), .B(SH[5]), .Y(n11) );
  NAND2BXL U356 ( .AN(SH[4]), .B(n75), .Y(n43) );
  NOR2BX1 U357 ( .AN(n12), .B(n3), .Y(B[8]) );
  NOR2XL U358 ( .A(n44), .B(SH[5]), .Y(n12) );
  NAND2BXL U359 ( .AN(SH[4]), .B(n76), .Y(n44) );
  NOR2BX1 U360 ( .AN(n13), .B(n3), .Y(B[9]) );
  NOR2XL U361 ( .A(n45), .B(SH[5]), .Y(n13) );
  NAND2BXL U362 ( .AN(SH[4]), .B(n77), .Y(n45) );
  NOR2BX1 U363 ( .AN(n14), .B(n3), .Y(B[10]) );
  NOR2XL U364 ( .A(n46), .B(SH[5]), .Y(n14) );
  NAND2BXL U365 ( .AN(SH[4]), .B(n78), .Y(n46) );
  NOR2BX1 U366 ( .AN(n15), .B(n3), .Y(B[11]) );
  NOR2XL U367 ( .A(n47), .B(SH[5]), .Y(n15) );
  NAND2BXL U368 ( .AN(SH[4]), .B(n79), .Y(n47) );
  NOR2BX1 U369 ( .AN(n16), .B(n3), .Y(B[12]) );
  NOR2XL U370 ( .A(n48), .B(SH[5]), .Y(n16) );
  NAND2BXL U371 ( .AN(SH[4]), .B(n80), .Y(n48) );
  NOR2BX1 U372 ( .AN(n17), .B(n3), .Y(B[13]) );
  NOR2XL U373 ( .A(n49), .B(SH[5]), .Y(n17) );
  NAND2BXL U374 ( .AN(SH[4]), .B(n81), .Y(n49) );
  NOR2BX1 U375 ( .AN(n18), .B(n3), .Y(B[14]) );
  NOR2XL U376 ( .A(n50), .B(SH[5]), .Y(n18) );
  NAND2BXL U377 ( .AN(SH[4]), .B(n82), .Y(n50) );
  NOR2BX1 U378 ( .AN(n19), .B(n3), .Y(B[15]) );
  NOR2XL U379 ( .A(n51), .B(SH[5]), .Y(n19) );
  NAND2BXL U380 ( .AN(SH[4]), .B(n83), .Y(n51) );
  NOR2BX1 U381 ( .AN(n20), .B(n3), .Y(B[16]) );
  NOR2XL U382 ( .A(n52), .B(SH[5]), .Y(n20) );
  MXI2XL U383 ( .A(n84), .B(n68), .S0(SH[4]), .Y(n52) );
  NOR2BX1 U384 ( .AN(n21), .B(n3), .Y(B[17]) );
  NOR2XL U385 ( .A(n53), .B(SH[5]), .Y(n21) );
  MXI2XL U386 ( .A(n85), .B(n69), .S0(SH[4]), .Y(n53) );
  NOR2BX1 U387 ( .AN(n22), .B(n3), .Y(B[18]) );
  NOR2XL U388 ( .A(n54), .B(SH[5]), .Y(n22) );
  MXI2XL U389 ( .A(n86), .B(n70), .S0(SH[4]), .Y(n54) );
  NOR2BX1 U390 ( .AN(n23), .B(n3), .Y(B[19]) );
  NOR2XL U391 ( .A(n55), .B(SH[5]), .Y(n23) );
  MXI2XL U392 ( .A(n87), .B(n71), .S0(SH[4]), .Y(n55) );
  NOR2BX1 U393 ( .AN(n24), .B(n3), .Y(B[20]) );
  NOR2XL U394 ( .A(n56), .B(SH[5]), .Y(n24) );
  MXI2XL U395 ( .A(n88), .B(n72), .S0(SH[4]), .Y(n56) );
  NOR2BX1 U396 ( .AN(n25), .B(n3), .Y(B[21]) );
  NOR2XL U397 ( .A(n57), .B(SH[5]), .Y(n25) );
  MXI2XL U398 ( .A(n89), .B(n73), .S0(SH[4]), .Y(n57) );
  NOR2BX1 U399 ( .AN(n26), .B(n3), .Y(B[22]) );
  NOR2XL U400 ( .A(n58), .B(SH[5]), .Y(n26) );
  MXI2XL U401 ( .A(n90), .B(n74), .S0(SH[4]), .Y(n58) );
  NOR2BX1 U402 ( .AN(n27), .B(n3), .Y(B[23]) );
  NOR2XL U403 ( .A(n59), .B(SH[5]), .Y(n27) );
  MXI2XL U404 ( .A(n91), .B(n75), .S0(SH[4]), .Y(n59) );
  NOR2BX1 U405 ( .AN(n28), .B(n3), .Y(B[24]) );
  NOR2XL U406 ( .A(n60), .B(SH[5]), .Y(n28) );
  MXI2XL U407 ( .A(n92), .B(n76), .S0(SH[4]), .Y(n60) );
  NOR2BX1 U408 ( .AN(n29), .B(n3), .Y(B[25]) );
  NOR2XL U409 ( .A(n61), .B(SH[5]), .Y(n29) );
  MXI2XL U410 ( .A(n93), .B(n77), .S0(SH[4]), .Y(n61) );
  NOR2BX1 U411 ( .AN(n30), .B(n3), .Y(B[26]) );
  NOR2XL U412 ( .A(n62), .B(SH[5]), .Y(n30) );
  MXI2XL U413 ( .A(n94), .B(n78), .S0(SH[4]), .Y(n62) );
  NOR2BX1 U414 ( .AN(n31), .B(n3), .Y(B[27]) );
  NOR2XL U415 ( .A(n63), .B(SH[5]), .Y(n31) );
  MXI2XL U416 ( .A(n95), .B(n79), .S0(SH[4]), .Y(n63) );
  NOR2BX1 U417 ( .AN(n32), .B(n3), .Y(B[28]) );
  NOR2XL U418 ( .A(n64), .B(SH[5]), .Y(n32) );
  MXI2XL U419 ( .A(n96), .B(n80), .S0(SH[4]), .Y(n64) );
  NOR2BX1 U420 ( .AN(n33), .B(n3), .Y(B[29]) );
  NOR2XL U421 ( .A(n65), .B(SH[5]), .Y(n33) );
  MXI2XL U422 ( .A(n97), .B(n81), .S0(SH[4]), .Y(n65) );
  NOR2BX1 U423 ( .AN(n34), .B(n3), .Y(B[30]) );
  NOR2XL U424 ( .A(n66), .B(SH[5]), .Y(n34) );
  MXI2XL U425 ( .A(n98), .B(n82), .S0(SH[4]), .Y(n66) );
  NOR2BX1 U426 ( .AN(n35), .B(n3), .Y(B[31]) );
  MXI2X1 U427 ( .A(n108), .B(n100), .S0(SH[3]), .Y(n76) );
  MXI2X1 U428 ( .A(n109), .B(n101), .S0(SH[3]), .Y(n77) );
  MXI2X1 U429 ( .A(n110), .B(n102), .S0(SH[3]), .Y(n78) );
  MXI2X1 U430 ( .A(n111), .B(n103), .S0(SH[3]), .Y(n79) );
  MXI2X1 U431 ( .A(n112), .B(n104), .S0(SH[3]), .Y(n80) );
  MXI2X1 U432 ( .A(n113), .B(n105), .S0(SH[3]), .Y(n81) );
  MXI2X1 U433 ( .A(n114), .B(n106), .S0(SH[3]), .Y(n82) );
  MXI2X1 U434 ( .A(n115), .B(n107), .S0(SH[3]), .Y(n83) );
  MXI2X1 U435 ( .A(n136), .B(n132), .S0(SH[2]), .Y(n104) );
  MXI2X1 U436 ( .A(n137), .B(n133), .S0(SH[2]), .Y(n105) );
  MXI2X1 U437 ( .A(n138), .B(n134), .S0(SH[2]), .Y(n106) );
  MXI2X1 U438 ( .A(n139), .B(n135), .S0(SH[2]), .Y(n107) );
  MXI2X1 U439 ( .A(n166), .B(n164), .S0(SH[1]), .Y(n134) );
  MXI2X1 U440 ( .A(n167), .B(n165), .S0(SH[1]), .Y(n135) );
  MXI2X1 U441 ( .A(n168), .B(n166), .S0(SH[1]), .Y(n136) );
  MXI2X1 U442 ( .A(n172), .B(n170), .S0(SH[1]), .Y(n140) );
  MXI2X1 U443 ( .A(n176), .B(n174), .S0(SH[1]), .Y(n144) );
  MXI2X1 U444 ( .A(n180), .B(n178), .S0(SH[1]), .Y(n148) );
  MXI2X1 U445 ( .A(n184), .B(n182), .S0(SH[1]), .Y(n152) );
  MXI2X1 U446 ( .A(n188), .B(n186), .S0(SH[1]), .Y(n156) );
  MXI2X1 U447 ( .A(n169), .B(n167), .S0(SH[1]), .Y(n137) );
  MXI2X1 U448 ( .A(n173), .B(n171), .S0(SH[1]), .Y(n141) );
  MXI2X1 U449 ( .A(n177), .B(n175), .S0(SH[1]), .Y(n145) );
  MXI2X1 U450 ( .A(n181), .B(n179), .S0(SH[1]), .Y(n149) );
  MXI2X1 U451 ( .A(n185), .B(n183), .S0(SH[1]), .Y(n153) );
  MXI2X1 U452 ( .A(n189), .B(n187), .S0(SH[1]), .Y(n157) );
  MXI2X1 U453 ( .A(n170), .B(n168), .S0(SH[1]), .Y(n138) );
  MXI2X1 U454 ( .A(n174), .B(n172), .S0(SH[1]), .Y(n142) );
  MXI2X1 U455 ( .A(n178), .B(n176), .S0(SH[1]), .Y(n146) );
  MXI2X1 U456 ( .A(n182), .B(n180), .S0(SH[1]), .Y(n150) );
  MXI2X1 U457 ( .A(n186), .B(n184), .S0(SH[1]), .Y(n154) );
  MXI2X1 U458 ( .A(n190), .B(n188), .S0(SH[1]), .Y(n158) );
  MXI2X1 U459 ( .A(n171), .B(n169), .S0(SH[1]), .Y(n139) );
  MXI2X1 U460 ( .A(n175), .B(n173), .S0(SH[1]), .Y(n143) );
  MXI2X1 U461 ( .A(n179), .B(n177), .S0(SH[1]), .Y(n147) );
  MXI2X1 U462 ( .A(n183), .B(n181), .S0(SH[1]), .Y(n151) );
  MXI2X1 U463 ( .A(n187), .B(n185), .S0(SH[1]), .Y(n155) );
  MXI2X1 U464 ( .A(n191), .B(n189), .S0(SH[1]), .Y(n159) );
  MXI2X1 U465 ( .A(n140), .B(n136), .S0(SH[2]), .Y(n108) );
  MXI2X1 U466 ( .A(n148), .B(n144), .S0(SH[2]), .Y(n116) );
  MXI2X1 U467 ( .A(n141), .B(n137), .S0(SH[2]), .Y(n109) );
  MXI2X1 U468 ( .A(n149), .B(n145), .S0(SH[2]), .Y(n117) );
  MXI2X1 U469 ( .A(n142), .B(n138), .S0(SH[2]), .Y(n110) );
  MXI2X1 U470 ( .A(n150), .B(n146), .S0(SH[2]), .Y(n118) );
  MXI2X1 U471 ( .A(n143), .B(n139), .S0(SH[2]), .Y(n111) );
  MXI2X1 U472 ( .A(n151), .B(n147), .S0(SH[2]), .Y(n119) );
  MXI2X1 U473 ( .A(n144), .B(n140), .S0(SH[2]), .Y(n112) );
  MXI2X1 U474 ( .A(n152), .B(n148), .S0(SH[2]), .Y(n120) );
  MXI2X1 U475 ( .A(n145), .B(n141), .S0(SH[2]), .Y(n113) );
  MXI2X1 U476 ( .A(n153), .B(n149), .S0(SH[2]), .Y(n121) );
  MXI2X1 U477 ( .A(n146), .B(n142), .S0(SH[2]), .Y(n114) );
  MXI2X1 U478 ( .A(n154), .B(n150), .S0(SH[2]), .Y(n122) );
  MXI2X1 U479 ( .A(n147), .B(n143), .S0(SH[2]), .Y(n115) );
  MXI2X1 U480 ( .A(n155), .B(n151), .S0(SH[2]), .Y(n123) );
  MXI2XL U481 ( .A(A[30]), .B(A[29]), .S0(SH[0]), .Y(n194) );
  MXI2XL U482 ( .A(A[31]), .B(A[30]), .S0(SH[0]), .Y(n195) );
  NOR2BX1 U483 ( .AN(n5), .B(n3), .Y(B[1]) );
  NOR2XL U484 ( .A(n37), .B(SH[5]), .Y(n5) );
  NAND2BXL U485 ( .AN(SH[4]), .B(n69), .Y(n37) );
  NAND2BXL U486 ( .AN(SH[0]), .B(A[0]), .Y(n164) );
  NAND2BXL U487 ( .AN(SH[2]), .B(n134), .Y(n102) );
  NAND2BXL U488 ( .AN(SH[2]), .B(n135), .Y(n103) );
  NAND2BXL U489 ( .AN(SH[2]), .B(n132), .Y(n100) );
  NAND2BXL U490 ( .AN(SH[2]), .B(n133), .Y(n101) );
  NAND2BXL U491 ( .AN(SH[4]), .B(n68), .Y(n36) );
  OR2X1 U492 ( .A(SH[15]), .B(SH[16]), .Y(n213) );
  OR2X1 U493 ( .A(SH[23]), .B(SH[24]), .Y(n217) );
  OR2X1 U494 ( .A(n205), .B(n204), .Y(n200) );
  OR2X1 U495 ( .A(n214), .B(n213), .Y(n205) );
  OR2X1 U496 ( .A(n216), .B(n215), .Y(n204) );
  OR2X1 U497 ( .A(SH[17]), .B(SH[18]), .Y(n214) );
  NAND2X1 U498 ( .A(n321), .B(n322), .Y(n207) );
  NAND2X1 U499 ( .A(n323), .B(n324), .Y(n202) );
  OR2X1 U500 ( .A(n203), .B(n208), .Y(n201) );
  OR2X1 U501 ( .A(n220), .B(n217), .Y(n203) );
  NAND2X1 U502 ( .A(n325), .B(n326), .Y(n206) );
  NOR2X1 U503 ( .A(SH[7]), .B(SH[6]), .Y(n326) );
endmodule


module alu_DW_rightsh_1 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n213, n214, n215,
         n216, n217, n220, n323, n324, n325, n326, n327, n328;

  MXI2XL U256 ( .A(A[30]), .B(A[31]), .S0(SH[0]), .Y(n194) );
  MXI2XL U257 ( .A(A[16]), .B(A[17]), .S0(SH[0]), .Y(n180) );
  MXI2XL U258 ( .A(A[6]), .B(A[7]), .S0(SH[0]), .Y(n170) );
  MXI2XL U259 ( .A(A[24]), .B(A[25]), .S0(SH[0]), .Y(n188) );
  MXI2XL U260 ( .A(A[17]), .B(A[18]), .S0(SH[0]), .Y(n181) );
  MXI2XL U261 ( .A(A[11]), .B(A[12]), .S0(SH[0]), .Y(n175) );
  MXI2XL U262 ( .A(A[25]), .B(A[26]), .S0(SH[0]), .Y(n189) );
  MXI2XL U263 ( .A(A[14]), .B(A[15]), .S0(SH[0]), .Y(n178) );
  MXI2XL U264 ( .A(A[15]), .B(A[16]), .S0(SH[0]), .Y(n179) );
  MXI2XL U265 ( .A(A[29]), .B(A[30]), .S0(SH[0]), .Y(n193) );
  MXI2XL U266 ( .A(A[4]), .B(A[5]), .S0(SH[0]), .Y(n168) );
  MXI2XL U267 ( .A(A[5]), .B(A[6]), .S0(SH[0]), .Y(n169) );
  MXI2XL U268 ( .A(A[22]), .B(A[23]), .S0(SH[0]), .Y(n186) );
  MXI2XL U269 ( .A(A[23]), .B(A[24]), .S0(SH[0]), .Y(n187) );
  MXI2XL U270 ( .A(A[18]), .B(A[19]), .S0(SH[0]), .Y(n182) );
  MXI2XL U271 ( .A(A[19]), .B(A[20]), .S0(SH[0]), .Y(n183) );
  MXI2XL U272 ( .A(A[20]), .B(A[21]), .S0(SH[0]), .Y(n184) );
  MXI2XL U273 ( .A(A[21]), .B(A[22]), .S0(SH[0]), .Y(n185) );
  MXI2XL U274 ( .A(A[12]), .B(A[13]), .S0(SH[0]), .Y(n176) );
  MXI2XL U275 ( .A(A[13]), .B(A[14]), .S0(SH[0]), .Y(n177) );
  MXI2XL U276 ( .A(A[9]), .B(A[10]), .S0(SH[0]), .Y(n173) );
  MXI2XL U277 ( .A(A[10]), .B(A[11]), .S0(SH[0]), .Y(n174) );
  MXI2XL U278 ( .A(A[2]), .B(A[3]), .S0(SH[0]), .Y(n166) );
  MXI2XL U279 ( .A(A[3]), .B(A[4]), .S0(SH[0]), .Y(n167) );
  MXI2XL U280 ( .A(A[7]), .B(A[8]), .S0(SH[0]), .Y(n171) );
  MXI2XL U281 ( .A(A[8]), .B(A[9]), .S0(SH[0]), .Y(n172) );
  MXI2XL U282 ( .A(A[26]), .B(A[27]), .S0(SH[0]), .Y(n190) );
  MXI2XL U283 ( .A(A[27]), .B(A[28]), .S0(SH[0]), .Y(n191) );
  MXI2XL U284 ( .A(n136), .B(n140), .S0(SH[2]), .Y(n104) );
  MXI2XL U285 ( .A(n137), .B(n141), .S0(SH[2]), .Y(n105) );
  MXI2XL U286 ( .A(n138), .B(n142), .S0(SH[2]), .Y(n106) );
  MXI2XL U287 ( .A(n139), .B(n143), .S0(SH[2]), .Y(n107) );
  NOR2XL U288 ( .A(n194), .B(SH[1]), .Y(n162) );
  NOR2XL U289 ( .A(n195), .B(SH[1]), .Y(n163) );
  NOR2XL U290 ( .A(n124), .B(SH[3]), .Y(n92) );
  NOR2XL U291 ( .A(n125), .B(SH[3]), .Y(n93) );
  NOR2XL U292 ( .A(n126), .B(SH[3]), .Y(n94) );
  NOR2XL U293 ( .A(n127), .B(SH[3]), .Y(n95) );
  NOR2XL U294 ( .A(n128), .B(SH[3]), .Y(n96) );
  NOR2XL U295 ( .A(n129), .B(SH[3]), .Y(n97) );
  NOR2XL U296 ( .A(n130), .B(SH[3]), .Y(n98) );
  NOR2XL U297 ( .A(n131), .B(SH[3]), .Y(n99) );
  MXI2XL U298 ( .A(n132), .B(n136), .S0(SH[2]), .Y(n100) );
  MXI2XL U299 ( .A(n164), .B(n166), .S0(SH[1]), .Y(n132) );
  MXI2XL U300 ( .A(n133), .B(n137), .S0(SH[2]), .Y(n101) );
  MXI2XL U301 ( .A(n165), .B(n167), .S0(SH[1]), .Y(n133) );
  MXI2XL U302 ( .A(n134), .B(n138), .S0(SH[2]), .Y(n102) );
  MXI2XL U303 ( .A(n166), .B(n168), .S0(SH[1]), .Y(n134) );
  MXI2XL U304 ( .A(n135), .B(n139), .S0(SH[2]), .Y(n103) );
  MXI2XL U305 ( .A(n167), .B(n169), .S0(SH[1]), .Y(n135) );
  MXI2XL U306 ( .A(n100), .B(n108), .S0(SH[3]), .Y(n68) );
  NOR2XL U307 ( .A(n37), .B(SH[5]), .Y(n5) );
  MXI2XL U308 ( .A(n69), .B(n85), .S0(SH[4]), .Y(n37) );
  MXI2XL U309 ( .A(n101), .B(n109), .S0(SH[3]), .Y(n69) );
  NOR2XL U310 ( .A(n38), .B(SH[5]), .Y(n6) );
  MXI2XL U311 ( .A(n70), .B(n86), .S0(SH[4]), .Y(n38) );
  MXI2XL U312 ( .A(n102), .B(n110), .S0(SH[3]), .Y(n70) );
  NOR2XL U313 ( .A(n39), .B(SH[5]), .Y(n7) );
  MXI2XL U314 ( .A(n71), .B(n87), .S0(SH[4]), .Y(n39) );
  MXI2XL U315 ( .A(n103), .B(n111), .S0(SH[3]), .Y(n71) );
  NOR2XL U316 ( .A(n40), .B(SH[5]), .Y(n8) );
  MXI2XL U317 ( .A(n72), .B(n88), .S0(SH[4]), .Y(n40) );
  MXI2XL U318 ( .A(n104), .B(n112), .S0(SH[3]), .Y(n72) );
  NOR2XL U319 ( .A(n41), .B(SH[5]), .Y(n9) );
  MXI2XL U320 ( .A(n73), .B(n89), .S0(SH[4]), .Y(n41) );
  MXI2XL U321 ( .A(n105), .B(n113), .S0(SH[3]), .Y(n73) );
  NOR2XL U322 ( .A(n42), .B(SH[5]), .Y(n10) );
  MXI2XL U323 ( .A(n74), .B(n90), .S0(SH[4]), .Y(n42) );
  MXI2XL U324 ( .A(n106), .B(n114), .S0(SH[3]), .Y(n74) );
  NOR2XL U325 ( .A(n43), .B(SH[5]), .Y(n11) );
  MXI2XL U326 ( .A(n75), .B(n91), .S0(SH[4]), .Y(n43) );
  MXI2XL U327 ( .A(n107), .B(n115), .S0(SH[3]), .Y(n75) );
  NOR2XL U328 ( .A(n44), .B(SH[5]), .Y(n12) );
  MXI2XL U329 ( .A(n76), .B(n92), .S0(SH[4]), .Y(n44) );
  MXI2XL U330 ( .A(n108), .B(n116), .S0(SH[3]), .Y(n76) );
  NOR2XL U331 ( .A(n45), .B(SH[5]), .Y(n13) );
  MXI2XL U332 ( .A(n77), .B(n93), .S0(SH[4]), .Y(n45) );
  MXI2XL U333 ( .A(n109), .B(n117), .S0(SH[3]), .Y(n77) );
  NOR2XL U334 ( .A(n46), .B(SH[5]), .Y(n14) );
  MXI2XL U335 ( .A(n78), .B(n94), .S0(SH[4]), .Y(n46) );
  MXI2XL U336 ( .A(n110), .B(n118), .S0(SH[3]), .Y(n78) );
  NOR2XL U337 ( .A(n52), .B(SH[5]), .Y(n20) );
  NOR2XL U338 ( .A(n53), .B(SH[5]), .Y(n21) );
  NOR2XL U339 ( .A(n54), .B(SH[5]), .Y(n22) );
  NOR2XL U340 ( .A(n55), .B(SH[5]), .Y(n23) );
  NOR2XL U341 ( .A(n56), .B(SH[5]), .Y(n24) );
  NOR2XL U342 ( .A(n57), .B(SH[5]), .Y(n25) );
  NOR2XL U343 ( .A(n58), .B(SH[5]), .Y(n26) );
  NOR2XL U344 ( .A(n59), .B(SH[5]), .Y(n27) );
  NOR2XL U345 ( .A(n60), .B(SH[5]), .Y(n28) );
  NOR2XL U346 ( .A(n61), .B(SH[5]), .Y(n29) );
  NOR2XL U347 ( .A(n62), .B(SH[5]), .Y(n30) );
  NOR2XL U348 ( .A(n63), .B(SH[5]), .Y(n31) );
  NOR2XL U349 ( .A(n64), .B(SH[5]), .Y(n32) );
  NOR2XL U350 ( .A(n65), .B(SH[5]), .Y(n33) );
  NOR2XL U351 ( .A(n66), .B(SH[5]), .Y(n34) );
  NOR2XL U352 ( .A(n67), .B(SH[5]), .Y(n35) );
  NOR2XL U353 ( .A(n47), .B(SH[5]), .Y(n15) );
  MXI2XL U354 ( .A(n79), .B(n95), .S0(SH[4]), .Y(n47) );
  MXI2XL U355 ( .A(n111), .B(n119), .S0(SH[3]), .Y(n79) );
  NOR2XL U356 ( .A(n48), .B(SH[5]), .Y(n16) );
  MXI2XL U357 ( .A(n80), .B(n96), .S0(SH[4]), .Y(n48) );
  MXI2XL U358 ( .A(n112), .B(n120), .S0(SH[3]), .Y(n80) );
  NOR2XL U359 ( .A(n49), .B(SH[5]), .Y(n17) );
  MXI2XL U360 ( .A(n81), .B(n97), .S0(SH[4]), .Y(n49) );
  MXI2XL U361 ( .A(n113), .B(n121), .S0(SH[3]), .Y(n81) );
  NOR2XL U362 ( .A(n50), .B(SH[5]), .Y(n18) );
  MXI2XL U363 ( .A(n82), .B(n98), .S0(SH[4]), .Y(n50) );
  MXI2XL U364 ( .A(n114), .B(n122), .S0(SH[3]), .Y(n82) );
  NOR2XL U365 ( .A(n51), .B(SH[5]), .Y(n19) );
  MXI2XL U366 ( .A(n83), .B(n99), .S0(SH[4]), .Y(n51) );
  MXI2XL U367 ( .A(n115), .B(n123), .S0(SH[3]), .Y(n83) );
  NOR2XL U368 ( .A(SH[9]), .B(SH[8]), .Y(n323) );
  NOR2XL U369 ( .A(SH[11]), .B(SH[10]), .Y(n324) );
  NOR2XL U370 ( .A(SH[25]), .B(SH[26]), .Y(n325) );
  NOR2XL U371 ( .A(SH[27]), .B(SH[28]), .Y(n326) );
  NOR2XL U372 ( .A(SH[13]), .B(SH[14]), .Y(n327) );
  OR2XL U373 ( .A(SH[19]), .B(SH[20]), .Y(n215) );
  OR2XL U374 ( .A(SH[21]), .B(SH[22]), .Y(n216) );
  OR2XL U375 ( .A(SH[31]), .B(SH[12]), .Y(n208) );
  OR2XL U376 ( .A(SH[29]), .B(SH[30]), .Y(n220) );
  OR2X6 U377 ( .A(n197), .B(n198), .Y(n3) );
  OR2X1 U378 ( .A(n199), .B(n200), .Y(n197) );
  OR2X1 U379 ( .A(n201), .B(n202), .Y(n198) );
  OR2X1 U380 ( .A(n206), .B(n207), .Y(n199) );
  MXI2X1 U381 ( .A(n116), .B(n124), .S0(SH[3]), .Y(n84) );
  MXI2X1 U382 ( .A(n117), .B(n125), .S0(SH[3]), .Y(n85) );
  MXI2X1 U383 ( .A(n118), .B(n126), .S0(SH[3]), .Y(n86) );
  MXI2X1 U384 ( .A(n119), .B(n127), .S0(SH[3]), .Y(n87) );
  MXI2X1 U385 ( .A(n120), .B(n128), .S0(SH[3]), .Y(n88) );
  MXI2X1 U386 ( .A(n121), .B(n129), .S0(SH[3]), .Y(n89) );
  MXI2X1 U387 ( .A(n122), .B(n130), .S0(SH[3]), .Y(n90) );
  MXI2X1 U388 ( .A(n123), .B(n131), .S0(SH[3]), .Y(n91) );
  MXI2X1 U389 ( .A(n156), .B(n160), .S0(SH[2]), .Y(n124) );
  MXI2X1 U390 ( .A(n157), .B(n161), .S0(SH[2]), .Y(n125) );
  MXI2X1 U391 ( .A(n158), .B(n162), .S0(SH[2]), .Y(n126) );
  MXI2X1 U392 ( .A(n159), .B(n163), .S0(SH[2]), .Y(n127) );
  MXI2X1 U393 ( .A(n192), .B(n194), .S0(SH[1]), .Y(n160) );
  MXI2X1 U394 ( .A(n193), .B(n195), .S0(SH[1]), .Y(n161) );
  MXI2X1 U395 ( .A(n168), .B(n170), .S0(SH[1]), .Y(n136) );
  MXI2X1 U396 ( .A(n169), .B(n171), .S0(SH[1]), .Y(n137) );
  MXI2X1 U397 ( .A(n170), .B(n172), .S0(SH[1]), .Y(n138) );
  MXI2X1 U398 ( .A(n171), .B(n173), .S0(SH[1]), .Y(n139) );
  MXI2X1 U399 ( .A(n172), .B(n174), .S0(SH[1]), .Y(n140) );
  MXI2X1 U400 ( .A(n173), .B(n175), .S0(SH[1]), .Y(n141) );
  MXI2X1 U401 ( .A(n174), .B(n176), .S0(SH[1]), .Y(n142) );
  MXI2X1 U402 ( .A(n175), .B(n177), .S0(SH[1]), .Y(n143) );
  MXI2X1 U403 ( .A(n176), .B(n178), .S0(SH[1]), .Y(n144) );
  MXI2X1 U404 ( .A(n177), .B(n179), .S0(SH[1]), .Y(n145) );
  MXI2X1 U405 ( .A(n178), .B(n180), .S0(SH[1]), .Y(n146) );
  MXI2X1 U406 ( .A(n179), .B(n181), .S0(SH[1]), .Y(n147) );
  MXI2X1 U407 ( .A(n180), .B(n182), .S0(SH[1]), .Y(n148) );
  MXI2X1 U408 ( .A(n181), .B(n183), .S0(SH[1]), .Y(n149) );
  MXI2X1 U409 ( .A(n182), .B(n184), .S0(SH[1]), .Y(n150) );
  MXI2X1 U410 ( .A(n183), .B(n185), .S0(SH[1]), .Y(n151) );
  MXI2X1 U411 ( .A(n184), .B(n186), .S0(SH[1]), .Y(n152) );
  MXI2X1 U412 ( .A(n185), .B(n187), .S0(SH[1]), .Y(n153) );
  MXI2X1 U413 ( .A(n186), .B(n188), .S0(SH[1]), .Y(n154) );
  MXI2X1 U414 ( .A(n187), .B(n189), .S0(SH[1]), .Y(n155) );
  MXI2X1 U415 ( .A(n188), .B(n190), .S0(SH[1]), .Y(n156) );
  MXI2X1 U416 ( .A(n189), .B(n191), .S0(SH[1]), .Y(n157) );
  MXI2X1 U417 ( .A(n190), .B(n192), .S0(SH[1]), .Y(n158) );
  MXI2X1 U418 ( .A(n191), .B(n193), .S0(SH[1]), .Y(n159) );
  MXI2XL U419 ( .A(A[28]), .B(A[29]), .S0(SH[0]), .Y(n192) );
  MXI2X1 U420 ( .A(n140), .B(n144), .S0(SH[2]), .Y(n108) );
  MXI2X1 U421 ( .A(n141), .B(n145), .S0(SH[2]), .Y(n109) );
  MXI2X1 U422 ( .A(n142), .B(n146), .S0(SH[2]), .Y(n110) );
  MXI2X1 U423 ( .A(n143), .B(n147), .S0(SH[2]), .Y(n111) );
  MXI2X1 U424 ( .A(n144), .B(n148), .S0(SH[2]), .Y(n112) );
  MXI2X1 U425 ( .A(n145), .B(n149), .S0(SH[2]), .Y(n113) );
  MXI2X1 U426 ( .A(n146), .B(n150), .S0(SH[2]), .Y(n114) );
  MXI2X1 U427 ( .A(n147), .B(n151), .S0(SH[2]), .Y(n115) );
  MXI2X1 U428 ( .A(n148), .B(n152), .S0(SH[2]), .Y(n116) );
  MXI2X1 U429 ( .A(n149), .B(n153), .S0(SH[2]), .Y(n117) );
  MXI2X1 U430 ( .A(n150), .B(n154), .S0(SH[2]), .Y(n118) );
  MXI2X1 U431 ( .A(n151), .B(n155), .S0(SH[2]), .Y(n119) );
  MXI2X1 U432 ( .A(n152), .B(n156), .S0(SH[2]), .Y(n120) );
  MXI2X1 U433 ( .A(n153), .B(n157), .S0(SH[2]), .Y(n121) );
  MXI2X1 U434 ( .A(n154), .B(n158), .S0(SH[2]), .Y(n122) );
  MXI2X1 U435 ( .A(n155), .B(n159), .S0(SH[2]), .Y(n123) );
  MXI2XL U436 ( .A(A[0]), .B(A[1]), .S0(SH[0]), .Y(n164) );
  MXI2XL U437 ( .A(A[1]), .B(A[2]), .S0(SH[0]), .Y(n165) );
  NAND2BXL U438 ( .AN(SH[0]), .B(A[31]), .Y(n195) );
  NAND2BXL U439 ( .AN(SH[2]), .B(n160), .Y(n128) );
  NAND2BXL U440 ( .AN(SH[2]), .B(n161), .Y(n129) );
  NAND2BXL U441 ( .AN(SH[2]), .B(n162), .Y(n130) );
  NAND2BXL U442 ( .AN(SH[2]), .B(n163), .Y(n131) );
  NOR2BX1 U443 ( .AN(n4), .B(n3), .Y(B[0]) );
  NOR2XL U444 ( .A(n36), .B(SH[5]), .Y(n4) );
  MXI2XL U445 ( .A(n68), .B(n84), .S0(SH[4]), .Y(n36) );
  NOR2BX1 U446 ( .AN(n5), .B(n3), .Y(B[1]) );
  NOR2BX1 U447 ( .AN(n6), .B(n3), .Y(B[2]) );
  NOR2BX1 U448 ( .AN(n7), .B(n3), .Y(B[3]) );
  NOR2BX1 U449 ( .AN(n8), .B(n3), .Y(B[4]) );
  NOR2BX1 U450 ( .AN(n9), .B(n3), .Y(B[5]) );
  NOR2BX1 U451 ( .AN(n10), .B(n3), .Y(B[6]) );
  NOR2BX1 U452 ( .AN(n11), .B(n3), .Y(B[7]) );
  NOR2BX1 U453 ( .AN(n12), .B(n3), .Y(B[8]) );
  NOR2BX1 U454 ( .AN(n13), .B(n3), .Y(B[9]) );
  NOR2BX1 U455 ( .AN(n14), .B(n3), .Y(B[10]) );
  NOR2BX1 U456 ( .AN(n15), .B(n3), .Y(B[11]) );
  NOR2BX1 U457 ( .AN(n16), .B(n3), .Y(B[12]) );
  NOR2BX1 U458 ( .AN(n17), .B(n3), .Y(B[13]) );
  NOR2BX1 U459 ( .AN(n18), .B(n3), .Y(B[14]) );
  NOR2BX1 U460 ( .AN(n19), .B(n3), .Y(B[15]) );
  NOR2BX1 U461 ( .AN(n20), .B(n3), .Y(B[16]) );
  NAND2BXL U462 ( .AN(SH[4]), .B(n84), .Y(n52) );
  NOR2BX1 U463 ( .AN(n21), .B(n3), .Y(B[17]) );
  NAND2BXL U464 ( .AN(SH[4]), .B(n85), .Y(n53) );
  NOR2BX1 U465 ( .AN(n22), .B(n3), .Y(B[18]) );
  NAND2BXL U466 ( .AN(SH[4]), .B(n86), .Y(n54) );
  NOR2BX1 U467 ( .AN(n23), .B(n3), .Y(B[19]) );
  NAND2BXL U468 ( .AN(SH[4]), .B(n87), .Y(n55) );
  NOR2BX1 U469 ( .AN(n24), .B(n3), .Y(B[20]) );
  NAND2BXL U470 ( .AN(SH[4]), .B(n88), .Y(n56) );
  NOR2BX1 U471 ( .AN(n25), .B(n3), .Y(B[21]) );
  NAND2BXL U472 ( .AN(SH[4]), .B(n89), .Y(n57) );
  NOR2BX1 U473 ( .AN(n26), .B(n3), .Y(B[22]) );
  NAND2BXL U474 ( .AN(SH[4]), .B(n90), .Y(n58) );
  NOR2BX1 U475 ( .AN(n27), .B(n3), .Y(B[23]) );
  NAND2BXL U476 ( .AN(SH[4]), .B(n91), .Y(n59) );
  NOR2BX1 U477 ( .AN(n28), .B(n3), .Y(B[24]) );
  NAND2BXL U478 ( .AN(SH[4]), .B(n92), .Y(n60) );
  NOR2BX1 U479 ( .AN(n29), .B(n3), .Y(B[25]) );
  NAND2BXL U480 ( .AN(SH[4]), .B(n93), .Y(n61) );
  NOR2BX1 U481 ( .AN(n30), .B(n3), .Y(B[26]) );
  NAND2BXL U482 ( .AN(SH[4]), .B(n94), .Y(n62) );
  NOR2BX1 U483 ( .AN(n31), .B(n3), .Y(B[27]) );
  NAND2BXL U484 ( .AN(SH[4]), .B(n95), .Y(n63) );
  NOR2BX1 U485 ( .AN(n32), .B(n3), .Y(B[28]) );
  NAND2BXL U486 ( .AN(SH[4]), .B(n96), .Y(n64) );
  NOR2BX1 U487 ( .AN(n33), .B(n3), .Y(B[29]) );
  NAND2BXL U488 ( .AN(SH[4]), .B(n97), .Y(n65) );
  NOR2BX1 U489 ( .AN(n34), .B(n3), .Y(B[30]) );
  NAND2BXL U490 ( .AN(SH[4]), .B(n98), .Y(n66) );
  NOR2BX1 U491 ( .AN(n35), .B(n3), .Y(B[31]) );
  NAND2BXL U492 ( .AN(SH[4]), .B(n99), .Y(n67) );
  OR2X1 U493 ( .A(SH[15]), .B(SH[16]), .Y(n213) );
  OR2X1 U494 ( .A(SH[23]), .B(SH[24]), .Y(n217) );
  OR2X1 U495 ( .A(n205), .B(n204), .Y(n200) );
  OR2X1 U496 ( .A(n214), .B(n213), .Y(n205) );
  OR2X1 U497 ( .A(n216), .B(n215), .Y(n204) );
  OR2X1 U498 ( .A(SH[17]), .B(SH[18]), .Y(n214) );
  NAND2X1 U499 ( .A(n323), .B(n324), .Y(n207) );
  NAND2X1 U500 ( .A(n325), .B(n326), .Y(n202) );
  OR2X1 U501 ( .A(n203), .B(n208), .Y(n201) );
  OR2X1 U502 ( .A(n220), .B(n217), .Y(n203) );
  NAND2X1 U503 ( .A(n327), .B(n328), .Y(n206) );
  NOR2X1 U504 ( .A(SH[7]), .B(SH[6]), .Y(n328) );
endmodule


module alu ( ALUin1, ALUin2, ALUctrl, ALUresult, ALUzero );
  input [31:0] ALUin1;
  input [31:0] ALUin2;
  input [3:0] ALUctrl;
  output [31:0] ALUresult;
  output ALUzero;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39,
         N40, N41, N42, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89,
         N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102,
         N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113,
         N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124,
         N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135,
         N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146,
         N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157,
         N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168,
         N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179,
         N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190,
         N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201,
         N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212,
         N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223,
         N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234,
         N235, N236, N237, N238, N271, N304, N305, N306, N307, N308, N309,
         N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331,
         N332, N333, N334, N335, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207;

  alu_DW01_addsub_0 r332 ( .A(ALUin1), .B(ALUin2), .CI(1'b0), .ADD_SUB(n2), 
        .SUM({N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, 
        N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, 
        N119, N118, N117, N116, N115, N114, N113, N112, N111}) );
  alu_DW01_cmp6_0 r323 ( .A(ALUin1), .B(ALUin2), .TC(1'b0), .LT(N271), .EQ(
        ALUzero) );
  alu_DW_leftsh_1 sll_1122 ( .A(ALUin1), .SH(ALUin2), .B({N174, N173, N172, 
        N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, 
        N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, 
        N147, N146, N145, N144, N143}) );
  alu_DW_rightsh_1 r321 ( .A(ALUin1), .DATA_TC(1'b0), .SH(ALUin2), .B({N206, 
        N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, 
        N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, 
        N181, N180, N179, N178, N177, N176, N175}) );
  AND2X2 U3 ( .A(N222), .B(n203), .Y(n99) );
  AND2X2 U6 ( .A(N221), .B(n203), .Y(n105) );
  AND2X2 U7 ( .A(N220), .B(n203), .Y(n111) );
  AND2X2 U8 ( .A(N216), .B(n203), .Y(n135) );
  AND2X2 U9 ( .A(N215), .B(n203), .Y(n141) );
  AND2X2 U10 ( .A(N214), .B(n203), .Y(n147) );
  AND2X2 U11 ( .A(N210), .B(n203), .Y(n171) );
  AND2X2 U12 ( .A(N209), .B(n203), .Y(n177) );
  AND2X2 U13 ( .A(N208), .B(n203), .Y(n183) );
  AND2X2 U14 ( .A(N207), .B(n203), .Y(n189) );
  AND2X2 U15 ( .A(N103), .B(n204), .Y(n46) );
  AND2X2 U16 ( .A(N231), .B(n203), .Y(n45) );
  AND2X2 U17 ( .A(N102), .B(n204), .Y(n52) );
  AND2X2 U18 ( .A(N230), .B(n203), .Y(n51) );
  AND2X2 U19 ( .A(N101), .B(n204), .Y(n58) );
  AND2X2 U20 ( .A(N229), .B(n203), .Y(n57) );
  AND2X2 U21 ( .A(N97), .B(n204), .Y(n82) );
  AND2X2 U22 ( .A(N225), .B(n203), .Y(n81) );
  AND2X2 U23 ( .A(N96), .B(n204), .Y(n88) );
  AND2X2 U24 ( .A(N224), .B(n203), .Y(n87) );
  AND2X2 U25 ( .A(N223), .B(n203), .Y(n93) );
  AND2X2 U26 ( .A(N219), .B(n203), .Y(n117) );
  AND2X2 U27 ( .A(N218), .B(n203), .Y(n123) );
  AND2X2 U28 ( .A(N217), .B(n203), .Y(n129) );
  AND2X2 U29 ( .A(N213), .B(n203), .Y(n153) );
  AND2X2 U30 ( .A(N212), .B(n203), .Y(n159) );
  AND2X2 U31 ( .A(N211), .B(n203), .Y(n165) );
  AND2X2 U32 ( .A(N100), .B(n204), .Y(n64) );
  AND2X2 U33 ( .A(N228), .B(n203), .Y(n63) );
  AND2X2 U34 ( .A(N99), .B(n204), .Y(n70) );
  AND2X2 U35 ( .A(N227), .B(n203), .Y(n69) );
  AND2X2 U36 ( .A(N98), .B(n204), .Y(n76) );
  AND2X2 U37 ( .A(N226), .B(n203), .Y(n75) );
  AND2X2 U38 ( .A(N107), .B(n204), .Y(n22) );
  AND2X2 U39 ( .A(N235), .B(n203), .Y(n21) );
  AND2X2 U40 ( .A(N108), .B(n204), .Y(n13) );
  AND2X2 U41 ( .A(N236), .B(n203), .Y(n12) );
  AND2X2 U42 ( .A(N106), .B(n204), .Y(n28) );
  AND2X2 U43 ( .A(N234), .B(n203), .Y(n27) );
  AND2X2 U44 ( .A(N105), .B(n204), .Y(n34) );
  AND2X2 U45 ( .A(N233), .B(n203), .Y(n33) );
  AND2X2 U46 ( .A(N104), .B(n204), .Y(n40) );
  NAND2X1 U47 ( .A(n203), .B(n204), .Y(n10) );
  AND2X2 U48 ( .A(N232), .B(n203), .Y(n39) );
  AND2X2 U49 ( .A(N109), .B(n204), .Y(n6) );
  AND2X2 U50 ( .A(N237), .B(n203), .Y(n5) );
  OAI211X1 U51 ( .A0(n204), .A1(n206), .B0(n201), .C0(n203), .Y(n9) );
  OR3X2 U52 ( .A(n207), .B(ALUctrl[3]), .C(ALUctrl[0]), .Y(n1) );
  INVX6 U53 ( .A(n1), .Y(n2) );
  NOR2XL U54 ( .A(ALUin2[0]), .B(ALUin1[0]), .Y(N238) );
  CLKBUFX6 U55 ( .A(n202), .Y(n3) );
  NAND2BXL U56 ( .AN(n11), .B(n3), .Y(n19) );
  NAND2BXL U57 ( .AN(n20), .B(n3), .Y(n25) );
  NAND2BXL U58 ( .AN(n26), .B(n3), .Y(n31) );
  NAND2BXL U59 ( .AN(n32), .B(n3), .Y(n37) );
  NAND2BXL U60 ( .AN(n38), .B(n3), .Y(n43) );
  NAND2BXL U61 ( .AN(n44), .B(n3), .Y(n49) );
  NAND2BXL U62 ( .AN(n50), .B(n3), .Y(n55) );
  NAND2BXL U63 ( .AN(n56), .B(n3), .Y(n61) );
  NAND2BXL U64 ( .AN(n62), .B(n3), .Y(n67) );
  NAND2BXL U65 ( .AN(n68), .B(n3), .Y(n73) );
  NAND2BXL U66 ( .AN(n74), .B(n3), .Y(n79) );
  NAND2BXL U67 ( .AN(n80), .B(n3), .Y(n85) );
  NAND2BXL U68 ( .AN(n86), .B(n3), .Y(n91) );
  NAND2BXL U69 ( .AN(n92), .B(n3), .Y(n97) );
  NAND2BXL U70 ( .AN(n98), .B(n3), .Y(n103) );
  NAND2BXL U71 ( .AN(n104), .B(n3), .Y(n109) );
  NAND2BXL U72 ( .AN(n110), .B(n3), .Y(n115) );
  NAND2BXL U73 ( .AN(n116), .B(n3), .Y(n121) );
  NAND2BXL U74 ( .AN(n122), .B(n3), .Y(n127) );
  NAND2BXL U75 ( .AN(n128), .B(n3), .Y(n133) );
  NAND2BXL U76 ( .AN(n134), .B(n3), .Y(n139) );
  NAND2BXL U77 ( .AN(n140), .B(n3), .Y(n145) );
  NAND2BXL U78 ( .AN(n146), .B(n3), .Y(n151) );
  NAND2BXL U79 ( .AN(n152), .B(n3), .Y(n157) );
  NAND2BXL U80 ( .AN(n158), .B(n3), .Y(n163) );
  NAND2BXL U81 ( .AN(n164), .B(n3), .Y(n169) );
  NAND2BXL U82 ( .AN(n170), .B(n3), .Y(n175) );
  NAND2BXL U83 ( .AN(n176), .B(n3), .Y(n181) );
  NAND2BXL U84 ( .AN(n182), .B(n3), .Y(n187) );
  NAND2BXL U85 ( .AN(n188), .B(n3), .Y(n193) );
  MXI2XL U86 ( .A(ALUctrl[3]), .B(n10), .S0(ALUctrl[0]), .Y(n202) );
  INVXL U87 ( .A(N237), .Y(N42) );
  INVXL U88 ( .A(N236), .Y(N41) );
  INVXL U89 ( .A(N235), .Y(N40) );
  XOR2XL U90 ( .A(ALUin2[27]), .B(ALUin1[27]), .Y(N308) );
  XOR2XL U91 ( .A(ALUin2[8]), .B(ALUin1[8]), .Y(N327) );
  XOR2XL U92 ( .A(ALUin2[26]), .B(ALUin1[26]), .Y(N309) );
  XOR2XL U93 ( .A(ALUin2[10]), .B(ALUin1[10]), .Y(N325) );
  XOR2XL U94 ( .A(ALUin2[3]), .B(ALUin1[3]), .Y(N332) );
  XOR2XL U95 ( .A(ALUin2[11]), .B(ALUin1[11]), .Y(N324) );
  XOR2XL U96 ( .A(ALUin2[13]), .B(ALUin1[13]), .Y(N322) );
  XOR2XL U97 ( .A(ALUin2[21]), .B(ALUin1[21]), .Y(N314) );
  XOR2XL U98 ( .A(ALUin2[12]), .B(ALUin1[12]), .Y(N323) );
  XOR2XL U99 ( .A(ALUin2[20]), .B(ALUin1[20]), .Y(N315) );
  XOR2XL U100 ( .A(ALUin2[9]), .B(ALUin1[9]), .Y(N326) );
  XOR2XL U101 ( .A(ALUin2[19]), .B(ALUin1[19]), .Y(N316) );
  XOR2XL U102 ( .A(ALUin2[22]), .B(ALUin1[22]), .Y(N313) );
  XOR2XL U103 ( .A(ALUin2[14]), .B(ALUin1[14]), .Y(N321) );
  XOR2XL U104 ( .A(ALUin2[28]), .B(ALUin1[28]), .Y(N307) );
  XOR2XL U105 ( .A(ALUin2[18]), .B(ALUin1[18]), .Y(N317) );
  XOR2XL U106 ( .A(ALUin2[2]), .B(ALUin1[2]), .Y(N333) );
  XOR2XL U107 ( .A(ALUin2[23]), .B(ALUin1[23]), .Y(N312) );
  XOR2XL U108 ( .A(ALUin2[5]), .B(ALUin1[5]), .Y(N330) );
  XOR2XL U109 ( .A(ALUin2[29]), .B(ALUin1[29]), .Y(N306) );
  XOR2XL U110 ( .A(ALUin2[15]), .B(ALUin1[15]), .Y(N320) );
  XOR2XL U111 ( .A(ALUin2[1]), .B(ALUin1[1]), .Y(N334) );
  XOR2XL U112 ( .A(ALUin2[24]), .B(ALUin1[24]), .Y(N311) );
  XOR2XL U113 ( .A(ALUin2[25]), .B(ALUin1[25]), .Y(N310) );
  XOR2XL U114 ( .A(ALUin2[4]), .B(ALUin1[4]), .Y(N331) );
  XOR2XL U115 ( .A(ALUin2[6]), .B(ALUin1[6]), .Y(N329) );
  XOR2XL U116 ( .A(ALUin2[7]), .B(ALUin1[7]), .Y(N328) );
  XOR2XL U117 ( .A(ALUin2[16]), .B(ALUin1[16]), .Y(N319) );
  XOR2XL U118 ( .A(ALUin2[17]), .B(ALUin1[17]), .Y(N318) );
  XOR2XL U119 ( .A(ALUin2[30]), .B(ALUin1[30]), .Y(N305) );
  XOR2XL U120 ( .A(ALUin2[31]), .B(ALUin1[31]), .Y(N304) );
  AND2XL U121 ( .A(ALUin2[0]), .B(ALUin1[0]), .Y(N110) );
  NAND2XL U122 ( .A(ALUctrl[2]), .B(ALUctrl[1]), .Y(n207) );
  NOR2XL U123 ( .A(ALUin2[1]), .B(ALUin1[1]), .Y(N237) );
  NOR2XL U124 ( .A(ALUin2[2]), .B(ALUin1[2]), .Y(N236) );
  NOR2XL U125 ( .A(ALUin2[3]), .B(ALUin1[3]), .Y(N235) );
  NOR2XL U126 ( .A(ALUin2[4]), .B(ALUin1[4]), .Y(N234) );
  NOR2XL U127 ( .A(ALUin2[5]), .B(ALUin1[5]), .Y(N233) );
  XNOR2XL U128 ( .A(ALUctrl[2]), .B(N238), .Y(n4) );
  NOR2XL U129 ( .A(ALUin2[9]), .B(ALUin1[9]), .Y(N229) );
  NOR2XL U130 ( .A(ALUin1[26]), .B(ALUin2[26]), .Y(N212) );
  NOR2XL U131 ( .A(ALUin2[19]), .B(ALUin1[19]), .Y(N219) );
  NOR2XL U132 ( .A(ALUin1[27]), .B(ALUin2[27]), .Y(N211) );
  NOR2XL U133 ( .A(ALUin2[10]), .B(ALUin1[10]), .Y(N228) );
  NOR2XL U134 ( .A(ALUin2[11]), .B(ALUin1[11]), .Y(N227) );
  NOR2XL U135 ( .A(ALUin2[13]), .B(ALUin1[13]), .Y(N225) );
  NOR2XL U136 ( .A(ALUin2[21]), .B(ALUin1[21]), .Y(N217) );
  NOR2XL U137 ( .A(ALUin2[12]), .B(ALUin1[12]), .Y(N226) );
  NOR2XL U138 ( .A(ALUin2[20]), .B(ALUin1[20]), .Y(N218) );
  NOR2XL U139 ( .A(ALUin2[8]), .B(ALUin1[8]), .Y(N230) );
  NOR2XL U140 ( .A(ALUin2[18]), .B(ALUin1[18]), .Y(N220) );
  NOR2XL U141 ( .A(ALUin2[14]), .B(ALUin1[14]), .Y(N224) );
  NOR2XL U142 ( .A(ALUin1[22]), .B(ALUin2[22]), .Y(N216) );
  NOR2XL U143 ( .A(ALUin1[28]), .B(ALUin2[28]), .Y(N210) );
  NOR2XL U144 ( .A(ALUin1[29]), .B(ALUin2[29]), .Y(N209) );
  NOR2XL U145 ( .A(ALUin2[15]), .B(ALUin1[15]), .Y(N223) );
  NOR2XL U146 ( .A(ALUin1[23]), .B(ALUin2[23]), .Y(N215) );
  NOR2XL U147 ( .A(ALUin2[6]), .B(ALUin1[6]), .Y(N232) );
  NOR2XL U148 ( .A(ALUin2[7]), .B(ALUin1[7]), .Y(N231) );
  NOR2XL U149 ( .A(ALUin2[16]), .B(ALUin1[16]), .Y(N222) );
  NOR2XL U150 ( .A(ALUin2[17]), .B(ALUin1[17]), .Y(N221) );
  NOR2XL U151 ( .A(ALUin1[24]), .B(ALUin2[24]), .Y(N214) );
  NOR2XL U152 ( .A(ALUin1[25]), .B(ALUin2[25]), .Y(N213) );
  NOR2XL U153 ( .A(ALUin1[30]), .B(ALUin2[30]), .Y(N208) );
  NOR2XL U154 ( .A(ALUin1[31]), .B(ALUin2[31]), .Y(N207) );
  AND2X2 U155 ( .A(N95), .B(n204), .Y(n94) );
  AND2X2 U156 ( .A(N94), .B(n204), .Y(n100) );
  MXI2X1 U157 ( .A(N111), .B(n195), .S0(ALUctrl[0]), .Y(n194) );
  MX2XL U158 ( .A(N143), .B(N271), .S0(ALUctrl[2]), .Y(n195) );
  MXI2X1 U159 ( .A(N175), .B(N335), .S0(ALUctrl[0]), .Y(n196) );
  MXI2X1 U160 ( .A(N113), .B(N145), .S0(ALUctrl[0]), .Y(n11) );
  MXI2X1 U161 ( .A(N114), .B(N146), .S0(ALUctrl[0]), .Y(n20) );
  MXI2X1 U162 ( .A(N115), .B(N147), .S0(ALUctrl[0]), .Y(n26) );
  MXI2X1 U163 ( .A(N116), .B(N148), .S0(ALUctrl[0]), .Y(n32) );
  MXI2X1 U164 ( .A(N117), .B(N149), .S0(ALUctrl[0]), .Y(n38) );
  MXI2X1 U165 ( .A(N118), .B(N150), .S0(ALUctrl[0]), .Y(n44) );
  MXI2X1 U166 ( .A(N119), .B(N151), .S0(ALUctrl[0]), .Y(n50) );
  MXI2X1 U167 ( .A(N120), .B(N152), .S0(ALUctrl[0]), .Y(n56) );
  MXI2X1 U168 ( .A(N121), .B(N153), .S0(ALUctrl[0]), .Y(n62) );
  MXI2X1 U169 ( .A(N122), .B(N154), .S0(ALUctrl[0]), .Y(n68) );
  MXI2X1 U170 ( .A(N123), .B(N155), .S0(ALUctrl[0]), .Y(n74) );
  MXI2X1 U171 ( .A(N124), .B(N156), .S0(ALUctrl[0]), .Y(n80) );
  MXI2X1 U172 ( .A(N125), .B(N157), .S0(ALUctrl[0]), .Y(n86) );
  MXI2X1 U173 ( .A(N126), .B(N158), .S0(ALUctrl[0]), .Y(n92) );
  MXI2X1 U174 ( .A(N127), .B(N159), .S0(ALUctrl[0]), .Y(n98) );
  MXI2X1 U175 ( .A(N128), .B(N160), .S0(ALUctrl[0]), .Y(n104) );
  MXI2X1 U176 ( .A(N129), .B(N161), .S0(ALUctrl[0]), .Y(n110) );
  MXI2X1 U177 ( .A(N130), .B(N162), .S0(ALUctrl[0]), .Y(n116) );
  MXI2X1 U178 ( .A(N131), .B(N163), .S0(ALUctrl[0]), .Y(n122) );
  MXI2X1 U179 ( .A(N132), .B(N164), .S0(ALUctrl[0]), .Y(n128) );
  MXI2X1 U180 ( .A(N133), .B(N165), .S0(ALUctrl[0]), .Y(n134) );
  MXI2X1 U181 ( .A(N134), .B(N166), .S0(ALUctrl[0]), .Y(n140) );
  MXI2X1 U182 ( .A(N135), .B(N167), .S0(ALUctrl[0]), .Y(n146) );
  MXI2X1 U183 ( .A(N136), .B(N168), .S0(ALUctrl[0]), .Y(n152) );
  MXI2X1 U184 ( .A(N137), .B(N169), .S0(ALUctrl[0]), .Y(n158) );
  MXI2X1 U185 ( .A(N138), .B(N170), .S0(ALUctrl[0]), .Y(n164) );
  MXI2X1 U186 ( .A(N139), .B(N171), .S0(ALUctrl[0]), .Y(n170) );
  MXI2X1 U187 ( .A(N140), .B(N172), .S0(ALUctrl[0]), .Y(n176) );
  MXI2X1 U188 ( .A(N141), .B(N173), .S0(ALUctrl[0]), .Y(n182) );
  MXI2X1 U189 ( .A(N142), .B(N174), .S0(ALUctrl[0]), .Y(n188) );
  INVX1 U190 ( .A(ALUctrl[0]), .Y(n206) );
  XOR2XL U191 ( .A(n204), .B(ALUctrl[3]), .Y(n200) );
  MX2XL U192 ( .A(N112), .B(N144), .S0(ALUctrl[0]), .Y(n201) );
  MX3XL U193 ( .A(n197), .B(n198), .C(n199), .S0(ALUctrl[3]), .S1(ALUctrl[1]), 
        .Y(ALUresult[0]) );
  NOR2BXL U194 ( .AN(n204), .B(n196), .Y(n198) );
  NOR2BXL U195 ( .AN(n203), .B(n194), .Y(n199) );
  MX3XL U196 ( .A(N110), .B(N175), .C(n4), .S0(ALUctrl[2]), .S1(ALUctrl[0]), 
        .Y(n197) );
  MXI3X1 U197 ( .A(n7), .B(n8), .C(n9), .S0(ALUctrl[0]), .S1(ALUctrl[1]), .Y(
        ALUresult[1]) );
  MXI3X1 U198 ( .A(N42), .B(N334), .C(n5), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n8) );
  MXI2X1 U199 ( .A(n6), .B(N176), .S0(n205), .Y(n7) );
  MXI3X1 U200 ( .A(n17), .B(n18), .C(n19), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[2]) );
  MXI3X1 U201 ( .A(N41), .B(N333), .C(n12), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n18) );
  MXI2X1 U202 ( .A(n13), .B(N177), .S0(n205), .Y(n17) );
  MXI3X1 U203 ( .A(n23), .B(n24), .C(n25), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[3]) );
  MXI3X1 U204 ( .A(N40), .B(N332), .C(n21), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n24) );
  MXI2X1 U205 ( .A(n22), .B(N178), .S0(n205), .Y(n23) );
  MXI3X1 U206 ( .A(n29), .B(n30), .C(n31), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[4]) );
  MXI3X1 U207 ( .A(N39), .B(N331), .C(n27), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n30) );
  MXI2X1 U208 ( .A(n28), .B(N179), .S0(n205), .Y(n29) );
  MXI3X1 U209 ( .A(n35), .B(n36), .C(n37), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[5]) );
  MXI3X1 U210 ( .A(N38), .B(N330), .C(n33), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n36) );
  MXI2X1 U211 ( .A(n34), .B(N180), .S0(n205), .Y(n35) );
  MXI3X1 U212 ( .A(n41), .B(n42), .C(n43), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[6]) );
  MXI3X1 U213 ( .A(N37), .B(N329), .C(n39), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n42) );
  MXI2X1 U214 ( .A(n40), .B(N181), .S0(n205), .Y(n41) );
  MXI3X1 U215 ( .A(n47), .B(n48), .C(n49), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[7]) );
  MXI3X1 U216 ( .A(N36), .B(N328), .C(n45), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n48) );
  MXI2X1 U217 ( .A(n46), .B(N182), .S0(n205), .Y(n47) );
  MXI3X1 U218 ( .A(n53), .B(n54), .C(n55), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[8]) );
  MXI3X1 U219 ( .A(N35), .B(N327), .C(n51), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n54) );
  MXI2X1 U220 ( .A(n52), .B(N183), .S0(n205), .Y(n53) );
  MXI3X1 U221 ( .A(n59), .B(n60), .C(n61), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[9]) );
  MXI3X1 U222 ( .A(N34), .B(N326), .C(n57), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n60) );
  MXI2X1 U223 ( .A(n58), .B(N184), .S0(n205), .Y(n59) );
  MXI3X1 U224 ( .A(n65), .B(n66), .C(n67), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[10]) );
  MXI3X1 U225 ( .A(N33), .B(N325), .C(n63), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n66) );
  MXI2X1 U226 ( .A(n64), .B(N185), .S0(n205), .Y(n65) );
  MXI3X1 U227 ( .A(n71), .B(n72), .C(n73), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[11]) );
  MXI3X1 U228 ( .A(N32), .B(N324), .C(n69), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n72) );
  MXI2XL U229 ( .A(n70), .B(N186), .S0(n205), .Y(n71) );
  MXI3X1 U230 ( .A(n77), .B(n78), .C(n79), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[12]) );
  MXI3X1 U231 ( .A(N31), .B(N323), .C(n75), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n78) );
  MXI2XL U232 ( .A(n76), .B(N187), .S0(n205), .Y(n77) );
  MXI3X1 U233 ( .A(n83), .B(n84), .C(n85), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[13]) );
  MXI3X1 U234 ( .A(N30), .B(N322), .C(n81), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n84) );
  MXI2XL U235 ( .A(n82), .B(N188), .S0(n205), .Y(n83) );
  MXI3X1 U236 ( .A(n89), .B(n90), .C(n91), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[14]) );
  MXI3X1 U237 ( .A(N29), .B(N321), .C(n87), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n90) );
  MXI2XL U238 ( .A(n88), .B(N189), .S0(n205), .Y(n89) );
  MXI3X1 U239 ( .A(n95), .B(n96), .C(n97), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[15]) );
  MXI3X1 U240 ( .A(N28), .B(N320), .C(n93), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n96) );
  MXI2XL U241 ( .A(n94), .B(N190), .S0(n205), .Y(n95) );
  MXI3X1 U242 ( .A(n101), .B(n102), .C(n103), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[16]) );
  MXI3X1 U243 ( .A(N27), .B(N319), .C(n99), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n102) );
  MXI2XL U244 ( .A(n100), .B(N191), .S0(n205), .Y(n101) );
  MXI3X1 U245 ( .A(n107), .B(n108), .C(n109), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[17]) );
  MXI3X1 U246 ( .A(N26), .B(N318), .C(n105), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n108) );
  MXI2XL U247 ( .A(n106), .B(N192), .S0(n205), .Y(n107) );
  MXI3X1 U248 ( .A(n113), .B(n114), .C(n115), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[18]) );
  MXI3X1 U249 ( .A(N25), .B(N317), .C(n111), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n114) );
  MXI2XL U250 ( .A(n112), .B(N193), .S0(n205), .Y(n113) );
  MXI3X1 U251 ( .A(n119), .B(n120), .C(n121), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[19]) );
  MXI3X1 U252 ( .A(N24), .B(N316), .C(n117), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n120) );
  MXI2XL U253 ( .A(n118), .B(N194), .S0(n205), .Y(n119) );
  MXI3X1 U254 ( .A(n125), .B(n126), .C(n127), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[20]) );
  MXI3X1 U255 ( .A(N23), .B(N315), .C(n123), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n126) );
  MXI2XL U256 ( .A(n124), .B(N195), .S0(n205), .Y(n125) );
  MXI3X1 U257 ( .A(n131), .B(n132), .C(n133), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[21]) );
  MXI3X1 U258 ( .A(N22), .B(N314), .C(n129), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n132) );
  MXI2XL U259 ( .A(n130), .B(N196), .S0(n205), .Y(n131) );
  MXI3X1 U260 ( .A(n137), .B(n138), .C(n139), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[22]) );
  MXI3X1 U261 ( .A(N21), .B(N313), .C(n135), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n138) );
  MXI2XL U262 ( .A(n136), .B(N197), .S0(n205), .Y(n137) );
  MXI3X1 U263 ( .A(n143), .B(n144), .C(n145), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[23]) );
  MXI3X1 U264 ( .A(N20), .B(N312), .C(n141), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n144) );
  MXI2XL U265 ( .A(n142), .B(N198), .S0(n205), .Y(n143) );
  MXI3X1 U266 ( .A(n149), .B(n150), .C(n151), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[24]) );
  MXI3X1 U267 ( .A(N19), .B(N311), .C(n147), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n150) );
  MXI2XL U268 ( .A(n148), .B(N199), .S0(n205), .Y(n149) );
  MXI3X1 U269 ( .A(n155), .B(n156), .C(n157), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[25]) );
  MXI3X1 U270 ( .A(N18), .B(N310), .C(n153), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n156) );
  MXI2XL U271 ( .A(n154), .B(N200), .S0(n205), .Y(n155) );
  MXI3X1 U272 ( .A(n161), .B(n162), .C(n163), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[26]) );
  MXI3X1 U273 ( .A(N17), .B(N309), .C(n159), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n162) );
  MXI2XL U274 ( .A(n160), .B(N201), .S0(n205), .Y(n161) );
  MXI3X1 U275 ( .A(n167), .B(n168), .C(n169), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[27]) );
  MXI3X1 U276 ( .A(N16), .B(N308), .C(n165), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n168) );
  MXI2XL U277 ( .A(n166), .B(N202), .S0(n205), .Y(n167) );
  MXI3X1 U278 ( .A(n173), .B(n174), .C(n175), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[28]) );
  MXI3X1 U279 ( .A(N15), .B(N307), .C(n171), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n174) );
  MXI2XL U280 ( .A(n172), .B(N203), .S0(n205), .Y(n173) );
  MXI3X1 U281 ( .A(n179), .B(n180), .C(n181), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[29]) );
  MXI3X1 U282 ( .A(N14), .B(N306), .C(n177), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n180) );
  MXI2XL U283 ( .A(n178), .B(N204), .S0(n205), .Y(n179) );
  MXI3X1 U284 ( .A(n185), .B(n186), .C(n187), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[30]) );
  MXI3X1 U285 ( .A(N13), .B(N305), .C(n183), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n186) );
  MXI2XL U286 ( .A(n184), .B(N205), .S0(n205), .Y(n185) );
  MXI3X1 U287 ( .A(n191), .B(n192), .C(n193), .S0(ALUctrl[0]), .S1(ALUctrl[1]), 
        .Y(ALUresult[31]) );
  MXI3X1 U288 ( .A(N12), .B(N304), .C(n189), .S0(ALUctrl[3]), .S1(ALUctrl[2]), 
        .Y(n192) );
  MXI2XL U289 ( .A(n190), .B(N206), .S0(n205), .Y(n191) );
  AND2X2 U290 ( .A(N93), .B(n204), .Y(n106) );
  AND2X2 U291 ( .A(N92), .B(n204), .Y(n112) );
  AND2X2 U292 ( .A(N91), .B(n204), .Y(n118) );
  AND2X2 U293 ( .A(N90), .B(n204), .Y(n124) );
  AND2X2 U294 ( .A(N89), .B(n204), .Y(n130) );
  AND2X2 U295 ( .A(N88), .B(n204), .Y(n136) );
  AND2X2 U296 ( .A(N87), .B(n204), .Y(n142) );
  AND2X2 U297 ( .A(N86), .B(n204), .Y(n148) );
  AND2X2 U298 ( .A(N85), .B(n204), .Y(n154) );
  AND2X2 U299 ( .A(N84), .B(n204), .Y(n160) );
  AND2X2 U300 ( .A(N83), .B(n204), .Y(n166) );
  AND2X2 U301 ( .A(N82), .B(n204), .Y(n172) );
  AND2XL U302 ( .A(N81), .B(n204), .Y(n178) );
  AND2XL U303 ( .A(N80), .B(n204), .Y(n184) );
  AND2XL U304 ( .A(N79), .B(n204), .Y(n190) );
  CLKINVX6 U305 ( .A(ALUctrl[3]), .Y(n203) );
  CLKINVX6 U306 ( .A(ALUctrl[2]), .Y(n204) );
  CLKINVX6 U307 ( .A(n200), .Y(n205) );
  AND2X1 U308 ( .A(ALUin1[11]), .B(ALUin2[11]), .Y(N99) );
  AND2X1 U309 ( .A(ALUin1[12]), .B(ALUin2[12]), .Y(N98) );
  AND2X1 U310 ( .A(ALUin1[13]), .B(ALUin2[13]), .Y(N97) );
  AND2X1 U311 ( .A(ALUin1[14]), .B(ALUin2[14]), .Y(N96) );
  AND2X1 U312 ( .A(ALUin1[15]), .B(ALUin2[15]), .Y(N95) );
  AND2X1 U313 ( .A(ALUin1[16]), .B(ALUin2[16]), .Y(N94) );
  AND2X1 U314 ( .A(ALUin1[17]), .B(ALUin2[17]), .Y(N93) );
  AND2X1 U315 ( .A(ALUin1[18]), .B(ALUin2[18]), .Y(N92) );
  AND2X1 U316 ( .A(ALUin1[19]), .B(ALUin2[19]), .Y(N91) );
  AND2X1 U317 ( .A(ALUin1[20]), .B(ALUin2[20]), .Y(N90) );
  AND2X1 U318 ( .A(ALUin1[21]), .B(ALUin2[21]), .Y(N89) );
  AND2X1 U319 ( .A(ALUin1[22]), .B(ALUin2[22]), .Y(N88) );
  AND2X1 U320 ( .A(ALUin1[23]), .B(ALUin2[23]), .Y(N87) );
  AND2X1 U321 ( .A(ALUin1[24]), .B(ALUin2[24]), .Y(N86) );
  AND2X1 U322 ( .A(ALUin1[25]), .B(ALUin2[25]), .Y(N85) );
  AND2X1 U323 ( .A(ALUin1[26]), .B(ALUin2[26]), .Y(N84) );
  AND2X1 U324 ( .A(ALUin1[27]), .B(ALUin2[27]), .Y(N83) );
  AND2X1 U325 ( .A(ALUin1[28]), .B(ALUin2[28]), .Y(N82) );
  AND2X1 U326 ( .A(ALUin1[29]), .B(ALUin2[29]), .Y(N81) );
  AND2X1 U327 ( .A(ALUin1[30]), .B(ALUin2[30]), .Y(N80) );
  AND2X1 U328 ( .A(ALUin1[31]), .B(ALUin2[31]), .Y(N79) );
  CLKINVX1 U329 ( .A(N234), .Y(N39) );
  CLKINVX1 U330 ( .A(N233), .Y(N38) );
  CLKINVX1 U331 ( .A(N232), .Y(N37) );
  CLKINVX1 U332 ( .A(N231), .Y(N36) );
  CLKINVX1 U333 ( .A(N230), .Y(N35) );
  CLKINVX1 U334 ( .A(N229), .Y(N34) );
  XOR2X1 U335 ( .A(ALUin2[0]), .B(ALUin1[0]), .Y(N335) );
  CLKINVX1 U336 ( .A(N228), .Y(N33) );
  CLKINVX1 U337 ( .A(N227), .Y(N32) );
  CLKINVX1 U338 ( .A(N226), .Y(N31) );
  CLKINVX1 U339 ( .A(N225), .Y(N30) );
  CLKINVX1 U340 ( .A(N224), .Y(N29) );
  CLKINVX1 U341 ( .A(N223), .Y(N28) );
  CLKINVX1 U342 ( .A(N222), .Y(N27) );
  CLKINVX1 U343 ( .A(N221), .Y(N26) );
  CLKINVX1 U344 ( .A(N220), .Y(N25) );
  CLKINVX1 U345 ( .A(N219), .Y(N24) );
  CLKINVX1 U346 ( .A(N218), .Y(N23) );
  CLKINVX1 U347 ( .A(N217), .Y(N22) );
  CLKINVX1 U348 ( .A(N216), .Y(N21) );
  CLKINVX1 U349 ( .A(N215), .Y(N20) );
  CLKINVX1 U350 ( .A(N214), .Y(N19) );
  CLKINVX1 U351 ( .A(N213), .Y(N18) );
  CLKINVX1 U352 ( .A(N212), .Y(N17) );
  CLKINVX1 U353 ( .A(N211), .Y(N16) );
  CLKINVX1 U354 ( .A(N210), .Y(N15) );
  CLKINVX1 U355 ( .A(N209), .Y(N14) );
  CLKINVX1 U356 ( .A(N208), .Y(N13) );
  CLKINVX1 U357 ( .A(N207), .Y(N12) );
  AND2X1 U358 ( .A(ALUin2[1]), .B(ALUin1[1]), .Y(N109) );
  AND2X1 U359 ( .A(ALUin2[2]), .B(ALUin1[2]), .Y(N108) );
  AND2X1 U360 ( .A(ALUin2[3]), .B(ALUin1[3]), .Y(N107) );
  AND2X1 U361 ( .A(ALUin2[4]), .B(ALUin1[4]), .Y(N106) );
  AND2X1 U362 ( .A(ALUin2[5]), .B(ALUin1[5]), .Y(N105) );
  AND2X1 U363 ( .A(ALUin2[6]), .B(ALUin1[6]), .Y(N104) );
  AND2X1 U364 ( .A(ALUin2[7]), .B(ALUin1[7]), .Y(N103) );
  AND2X1 U365 ( .A(ALUin2[8]), .B(ALUin1[8]), .Y(N102) );
  AND2X1 U366 ( .A(ALUin2[9]), .B(ALUin1[9]), .Y(N101) );
  AND2X1 U367 ( .A(ALUin2[10]), .B(ALUin1[10]), .Y(N100) );
endmodule


module EXMEM ( clk, WB, M, ALUOut, RegRD, writedata, EX_pcplus4, WB_reg, M_reg, 
        ALUOut_reg, RegRD_reg, Writedata_reg, stall_bothzero, MEM_pcplus4 );
  input [2:0] WB;
  input [2:0] M;
  input [31:0] ALUOut;
  input [4:0] RegRD;
  input [31:0] writedata;
  input [31:0] EX_pcplus4;
  output [2:0] WB_reg;
  output [2:0] M_reg;
  output [31:0] ALUOut_reg;
  output [4:0] RegRD_reg;
  output [31:0] Writedata_reg;
  output [31:0] MEM_pcplus4;
  input clk, stall_bothzero;
  wire   n127, n128, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n117, n119, n120, n121, n122, n123, n124, n125, n126;

  EDFFX1 \WB_reg_reg[0]  ( .D(WB[0]), .E(n124), .CK(clk), .Q(WB_reg[0]) );
  EDFFX1 \ALUOut_reg_reg[1]  ( .D(ALUOut[1]), .E(stall_bothzero), .CK(clk), 
        .Q(ALUOut_reg[1]) );
  EDFFX1 \ALUOut_reg_reg[0]  ( .D(ALUOut[0]), .E(n126), .CK(clk), .Q(
        ALUOut_reg[0]) );
  EDFFX1 \RegRD_reg_reg[2]  ( .D(RegRD[2]), .E(n123), .CK(clk), .Q(
        RegRD_reg[2]) );
  EDFFX1 \RegRD_reg_reg[3]  ( .D(RegRD[3]), .E(n123), .CK(clk), .Q(
        RegRD_reg[3]) );
  EDFFX1 \RegRD_reg_reg[4]  ( .D(RegRD[4]), .E(n123), .CK(clk), .Q(
        RegRD_reg[4]) );
  EDFFX1 \RegRD_reg_reg[0]  ( .D(RegRD[0]), .E(n123), .CK(clk), .Q(
        RegRD_reg[0]) );
  EDFFX1 \RegRD_reg_reg[1]  ( .D(RegRD[1]), .E(n123), .CK(clk), .Q(
        RegRD_reg[1]) );
  EDFFX1 \ALUOut_reg_reg[6]  ( .D(ALUOut[6]), .E(n125), .CK(clk), .Q(
        ALUOut_reg[6]) );
  EDFFX1 \ALUOut_reg_reg[5]  ( .D(ALUOut[5]), .E(n125), .CK(clk), .Q(
        ALUOut_reg[5]) );
  EDFFX1 \ALUOut_reg_reg[4]  ( .D(ALUOut[4]), .E(n124), .CK(clk), .Q(
        ALUOut_reg[4]) );
  EDFFX1 \M_reg_reg[2]  ( .D(M[2]), .E(n123), .CK(clk), .Q(M_reg[2]) );
  EDFFX1 \MEM_pcplus4_reg[31]  ( .D(EX_pcplus4[31]), .E(n119), .CK(clk), .Q(
        MEM_pcplus4[31]) );
  EDFFX1 \MEM_pcplus4_reg[30]  ( .D(EX_pcplus4[30]), .E(n119), .CK(clk), .Q(
        MEM_pcplus4[30]) );
  EDFFX1 \MEM_pcplus4_reg[29]  ( .D(EX_pcplus4[29]), .E(n119), .CK(clk), .Q(
        MEM_pcplus4[29]) );
  EDFFX1 \MEM_pcplus4_reg[28]  ( .D(EX_pcplus4[28]), .E(n119), .CK(clk), .Q(
        MEM_pcplus4[28]) );
  EDFFX1 \MEM_pcplus4_reg[27]  ( .D(EX_pcplus4[27]), .E(n119), .CK(clk), .Q(
        MEM_pcplus4[27]) );
  EDFFX1 \MEM_pcplus4_reg[26]  ( .D(EX_pcplus4[26]), .E(n119), .CK(clk), .Q(
        MEM_pcplus4[26]) );
  EDFFX1 \M_reg_reg[0]  ( .D(M[0]), .E(n123), .CK(clk), .Q(M_reg[0]) );
  EDFFX1 \MEM_pcplus4_reg[25]  ( .D(EX_pcplus4[25]), .E(n120), .CK(clk), .Q(
        MEM_pcplus4[25]) );
  EDFFX1 \MEM_pcplus4_reg[24]  ( .D(EX_pcplus4[24]), .E(n120), .CK(clk), .Q(
        MEM_pcplus4[24]) );
  EDFFX1 \MEM_pcplus4_reg[23]  ( .D(EX_pcplus4[23]), .E(n120), .CK(clk), .Q(
        MEM_pcplus4[23]) );
  EDFFX1 \MEM_pcplus4_reg[22]  ( .D(EX_pcplus4[22]), .E(n120), .CK(clk), .Q(
        MEM_pcplus4[22]) );
  EDFFX1 \MEM_pcplus4_reg[21]  ( .D(EX_pcplus4[21]), .E(n120), .CK(clk), .Q(
        MEM_pcplus4[21]) );
  EDFFX1 \MEM_pcplus4_reg[20]  ( .D(EX_pcplus4[20]), .E(n120), .CK(clk), .Q(
        MEM_pcplus4[20]) );
  EDFFX1 \MEM_pcplus4_reg[19]  ( .D(EX_pcplus4[19]), .E(n120), .CK(clk), .Q(
        MEM_pcplus4[19]) );
  EDFFX1 \MEM_pcplus4_reg[18]  ( .D(EX_pcplus4[18]), .E(n121), .CK(clk), .Q(
        MEM_pcplus4[18]) );
  EDFFX1 \MEM_pcplus4_reg[17]  ( .D(EX_pcplus4[17]), .E(n121), .CK(clk), .Q(
        MEM_pcplus4[17]) );
  EDFFX1 \MEM_pcplus4_reg[16]  ( .D(EX_pcplus4[16]), .E(n121), .CK(clk), .Q(
        MEM_pcplus4[16]) );
  EDFFX1 \MEM_pcplus4_reg[15]  ( .D(EX_pcplus4[15]), .E(n121), .CK(clk), .Q(
        MEM_pcplus4[15]) );
  EDFFX1 \MEM_pcplus4_reg[14]  ( .D(EX_pcplus4[14]), .E(n121), .CK(clk), .Q(
        MEM_pcplus4[14]) );
  EDFFX1 \MEM_pcplus4_reg[13]  ( .D(EX_pcplus4[13]), .E(n121), .CK(clk), .Q(
        MEM_pcplus4[13]) );
  EDFFX1 \MEM_pcplus4_reg[12]  ( .D(EX_pcplus4[12]), .E(n121), .CK(clk), .Q(
        MEM_pcplus4[12]) );
  EDFFX1 \MEM_pcplus4_reg[11]  ( .D(EX_pcplus4[11]), .E(n122), .CK(clk), .Q(
        MEM_pcplus4[11]) );
  EDFFX1 \MEM_pcplus4_reg[10]  ( .D(EX_pcplus4[10]), .E(n122), .CK(clk), .Q(
        MEM_pcplus4[10]) );
  EDFFX1 \MEM_pcplus4_reg[9]  ( .D(EX_pcplus4[9]), .E(n122), .CK(clk), .Q(
        MEM_pcplus4[9]) );
  EDFFX1 \MEM_pcplus4_reg[8]  ( .D(EX_pcplus4[8]), .E(n122), .CK(clk), .Q(
        MEM_pcplus4[8]) );
  EDFFX1 \MEM_pcplus4_reg[7]  ( .D(EX_pcplus4[7]), .E(n122), .CK(clk), .Q(
        MEM_pcplus4[7]) );
  EDFFX1 \MEM_pcplus4_reg[6]  ( .D(EX_pcplus4[6]), .E(n123), .CK(clk), .Q(
        MEM_pcplus4[6]) );
  EDFFX1 \MEM_pcplus4_reg[5]  ( .D(EX_pcplus4[5]), .E(n123), .CK(clk), .Q(
        MEM_pcplus4[5]) );
  EDFFX1 \MEM_pcplus4_reg[4]  ( .D(EX_pcplus4[4]), .E(n123), .CK(clk), .Q(
        MEM_pcplus4[4]) );
  EDFFX1 \MEM_pcplus4_reg[3]  ( .D(EX_pcplus4[3]), .E(n124), .CK(clk), .Q(
        MEM_pcplus4[3]) );
  EDFFX1 \MEM_pcplus4_reg[2]  ( .D(EX_pcplus4[2]), .E(n124), .CK(clk), .Q(
        MEM_pcplus4[2]) );
  EDFFX1 \MEM_pcplus4_reg[1]  ( .D(EX_pcplus4[1]), .E(n120), .CK(clk), .Q(
        MEM_pcplus4[1]) );
  EDFFX1 \MEM_pcplus4_reg[0]  ( .D(EX_pcplus4[0]), .E(stall_bothzero), .CK(clk), .Q(MEM_pcplus4[0]) );
  EDFFX1 \WB_reg_reg[2]  ( .D(WB[2]), .E(n124), .CK(clk), .Q(WB_reg[2]) );
  EDFFX1 \WB_reg_reg[1]  ( .D(WB[1]), .E(n123), .CK(clk), .Q(WB_reg[1]) );
  EDFFX1 \M_reg_reg[1]  ( .D(M[1]), .E(n124), .CK(clk), .QN(n117) );
  EDFFX1 \ALUOut_reg_reg[2]  ( .D(ALUOut[2]), .E(n126), .CK(clk), .Q(n128) );
  EDFFX1 \ALUOut_reg_reg[3]  ( .D(ALUOut[3]), .E(n124), .CK(clk), .Q(n127) );
  EDFFX1 \ALUOut_reg_reg[12]  ( .D(ALUOut[12]), .E(n124), .CK(clk), .QN(n13)
         );
  EDFFX1 \ALUOut_reg_reg[11]  ( .D(ALUOut[11]), .E(n124), .CK(clk), .QN(n14)
         );
  EDFFX1 \ALUOut_reg_reg[10]  ( .D(ALUOut[10]), .E(n125), .CK(clk), .QN(n15)
         );
  EDFFX1 \ALUOut_reg_reg[27]  ( .D(ALUOut[27]), .E(n125), .CK(clk), .QN(n5) );
  EDFFX1 \ALUOut_reg_reg[26]  ( .D(ALUOut[26]), .E(n126), .CK(clk), .QN(n6) );
  EDFFX1 \ALUOut_reg_reg[25]  ( .D(ALUOut[25]), .E(n126), .CK(clk), .QN(n7) );
  EDFFX1 \ALUOut_reg_reg[21]  ( .D(ALUOut[21]), .E(n125), .CK(clk), .QN(n8) );
  EDFFX1 \ALUOut_reg_reg[20]  ( .D(ALUOut[20]), .E(n125), .CK(clk), .QN(n9) );
  EDFFX1 \ALUOut_reg_reg[19]  ( .D(ALUOut[19]), .E(n125), .CK(clk), .QN(n10)
         );
  EDFFX1 \ALUOut_reg_reg[15]  ( .D(ALUOut[15]), .E(n125), .CK(clk), .QN(n11)
         );
  EDFFX1 \ALUOut_reg_reg[14]  ( .D(ALUOut[14]), .E(n126), .CK(clk), .QN(n12)
         );
  EDFFX1 \ALUOut_reg_reg[13]  ( .D(ALUOut[13]), .E(n126), .CK(clk), .QN(n1) );
  EDFFX1 \ALUOut_reg_reg[9]  ( .D(ALUOut[9]), .E(n126), .CK(clk), .QN(n2) );
  EDFFX1 \ALUOut_reg_reg[8]  ( .D(ALUOut[8]), .E(n126), .CK(clk), .QN(n3) );
  EDFFX1 \ALUOut_reg_reg[7]  ( .D(ALUOut[7]), .E(n125), .CK(clk), .QN(n4) );
  EDFFX1 \ALUOut_reg_reg[31]  ( .D(ALUOut[31]), .E(n126), .CK(clk), .QN(n16)
         );
  EDFFX1 \ALUOut_reg_reg[30]  ( .D(ALUOut[30]), .E(n126), .CK(clk), .QN(n17)
         );
  EDFFX1 \ALUOut_reg_reg[29]  ( .D(ALUOut[29]), .E(n125), .CK(clk), .QN(n18)
         );
  EDFFX1 \ALUOut_reg_reg[28]  ( .D(ALUOut[28]), .E(n125), .CK(clk), .QN(n19)
         );
  EDFFX1 \ALUOut_reg_reg[24]  ( .D(ALUOut[24]), .E(n125), .CK(clk), .QN(n20)
         );
  EDFFX1 \ALUOut_reg_reg[23]  ( .D(ALUOut[23]), .E(n125), .CK(clk), .QN(n21)
         );
  EDFFX1 \ALUOut_reg_reg[22]  ( .D(ALUOut[22]), .E(n126), .CK(clk), .QN(n22)
         );
  EDFFX1 \ALUOut_reg_reg[18]  ( .D(ALUOut[18]), .E(n124), .CK(clk), .QN(n23)
         );
  EDFFX1 \ALUOut_reg_reg[17]  ( .D(ALUOut[17]), .E(n126), .CK(clk), .QN(n24)
         );
  EDFFX1 \ALUOut_reg_reg[16]  ( .D(ALUOut[16]), .E(n126), .CK(clk), .QN(n25)
         );
  EDFFX1 \Writedata_reg_reg[31]  ( .D(writedata[31]), .E(n119), .CK(clk), .QN(
        n26) );
  EDFFX1 \Writedata_reg_reg[30]  ( .D(writedata[30]), .E(n119), .CK(clk), .QN(
        n27) );
  EDFFX1 \Writedata_reg_reg[29]  ( .D(writedata[29]), .E(n119), .CK(clk), .QN(
        n28) );
  EDFFX1 \Writedata_reg_reg[28]  ( .D(writedata[28]), .E(n119), .CK(clk), .QN(
        n29) );
  EDFFX1 \Writedata_reg_reg[27]  ( .D(writedata[27]), .E(n119), .CK(clk), .QN(
        n30) );
  EDFFX1 \Writedata_reg_reg[26]  ( .D(writedata[26]), .E(n119), .CK(clk), .QN(
        n31) );
  EDFFX1 \Writedata_reg_reg[25]  ( .D(writedata[25]), .E(n119), .CK(clk), .QN(
        n32) );
  EDFFX1 \Writedata_reg_reg[24]  ( .D(writedata[24]), .E(n120), .CK(clk), .QN(
        n33) );
  EDFFX1 \Writedata_reg_reg[23]  ( .D(writedata[23]), .E(n120), .CK(clk), .QN(
        n34) );
  EDFFX1 \Writedata_reg_reg[22]  ( .D(writedata[22]), .E(n120), .CK(clk), .QN(
        n35) );
  EDFFX1 \Writedata_reg_reg[21]  ( .D(writedata[21]), .E(n120), .CK(clk), .QN(
        n36) );
  EDFFX1 \Writedata_reg_reg[20]  ( .D(writedata[20]), .E(n120), .CK(clk), .QN(
        n37) );
  EDFFX1 \Writedata_reg_reg[19]  ( .D(writedata[19]), .E(n120), .CK(clk), .QN(
        n38) );
  EDFFX1 \Writedata_reg_reg[18]  ( .D(writedata[18]), .E(n124), .CK(clk), .QN(
        n39) );
  EDFFX1 \Writedata_reg_reg[17]  ( .D(writedata[17]), .E(n121), .CK(clk), .QN(
        n40) );
  EDFFX1 \Writedata_reg_reg[16]  ( .D(writedata[16]), .E(n121), .CK(clk), .QN(
        n41) );
  EDFFX1 \Writedata_reg_reg[15]  ( .D(writedata[15]), .E(n121), .CK(clk), .QN(
        n42) );
  EDFFX1 \Writedata_reg_reg[14]  ( .D(writedata[14]), .E(n121), .CK(clk), .QN(
        n43) );
  EDFFX1 \Writedata_reg_reg[13]  ( .D(writedata[13]), .E(n121), .CK(clk), .QN(
        n44) );
  EDFFX1 \Writedata_reg_reg[12]  ( .D(writedata[12]), .E(n121), .CK(clk), .QN(
        n45) );
  EDFFX1 \Writedata_reg_reg[11]  ( .D(writedata[11]), .E(n122), .CK(clk), .QN(
        n46) );
  EDFFX1 \Writedata_reg_reg[10]  ( .D(writedata[10]), .E(n122), .CK(clk), .QN(
        n47) );
  EDFFX1 \Writedata_reg_reg[9]  ( .D(writedata[9]), .E(n122), .CK(clk), .QN(
        n48) );
  EDFFX1 \Writedata_reg_reg[8]  ( .D(writedata[8]), .E(n122), .CK(clk), .QN(
        n49) );
  EDFFX1 \Writedata_reg_reg[7]  ( .D(writedata[7]), .E(n122), .CK(clk), .QN(
        n50) );
  EDFFX1 \Writedata_reg_reg[6]  ( .D(writedata[6]), .E(n122), .CK(clk), .QN(
        n51) );
  EDFFX1 \Writedata_reg_reg[5]  ( .D(writedata[5]), .E(n122), .CK(clk), .QN(
        n52) );
  EDFFX1 \Writedata_reg_reg[4]  ( .D(writedata[4]), .E(n124), .CK(clk), .QN(
        n53) );
  EDFFX1 \Writedata_reg_reg[3]  ( .D(writedata[3]), .E(n122), .CK(clk), .QN(
        n54) );
  EDFFX1 \Writedata_reg_reg[2]  ( .D(writedata[2]), .E(n123), .CK(clk), .QN(
        n55) );
  EDFFX1 \Writedata_reg_reg[1]  ( .D(writedata[1]), .E(n124), .CK(clk), .QN(
        n56) );
  EDFFX1 \Writedata_reg_reg[0]  ( .D(writedata[0]), .E(n123), .CK(clk), .QN(
        n57) );
  INVX16 U2 ( .A(n57), .Y(Writedata_reg[0]) );
  INVX16 U3 ( .A(n56), .Y(Writedata_reg[1]) );
  INVX16 U4 ( .A(n55), .Y(Writedata_reg[2]) );
  INVX16 U5 ( .A(n54), .Y(Writedata_reg[3]) );
  INVX16 U6 ( .A(n53), .Y(Writedata_reg[4]) );
  INVX16 U7 ( .A(n52), .Y(Writedata_reg[5]) );
  INVX16 U8 ( .A(n51), .Y(Writedata_reg[6]) );
  INVX16 U9 ( .A(n50), .Y(Writedata_reg[7]) );
  INVX16 U10 ( .A(n49), .Y(Writedata_reg[8]) );
  INVX16 U11 ( .A(n48), .Y(Writedata_reg[9]) );
  INVX16 U12 ( .A(n47), .Y(Writedata_reg[10]) );
  INVX16 U13 ( .A(n46), .Y(Writedata_reg[11]) );
  INVX16 U14 ( .A(n45), .Y(Writedata_reg[12]) );
  INVX16 U15 ( .A(n44), .Y(Writedata_reg[13]) );
  INVX16 U16 ( .A(n43), .Y(Writedata_reg[14]) );
  INVX16 U17 ( .A(n42), .Y(Writedata_reg[15]) );
  INVX16 U18 ( .A(n41), .Y(Writedata_reg[16]) );
  INVX16 U19 ( .A(n40), .Y(Writedata_reg[17]) );
  INVX16 U20 ( .A(n39), .Y(Writedata_reg[18]) );
  INVX16 U21 ( .A(n38), .Y(Writedata_reg[19]) );
  INVX16 U22 ( .A(n37), .Y(Writedata_reg[20]) );
  INVX16 U23 ( .A(n36), .Y(Writedata_reg[21]) );
  INVX16 U24 ( .A(n35), .Y(Writedata_reg[22]) );
  INVX16 U25 ( .A(n34), .Y(Writedata_reg[23]) );
  INVX16 U26 ( .A(n33), .Y(Writedata_reg[24]) );
  INVX16 U27 ( .A(n32), .Y(Writedata_reg[25]) );
  INVX16 U28 ( .A(n31), .Y(Writedata_reg[26]) );
  INVX16 U29 ( .A(n30), .Y(Writedata_reg[27]) );
  INVX16 U30 ( .A(n29), .Y(Writedata_reg[28]) );
  INVX16 U31 ( .A(n28), .Y(Writedata_reg[29]) );
  INVX16 U32 ( .A(n27), .Y(Writedata_reg[30]) );
  INVX16 U33 ( .A(n26), .Y(Writedata_reg[31]) );
  INVX16 U34 ( .A(n25), .Y(ALUOut_reg[16]) );
  INVX16 U35 ( .A(n24), .Y(ALUOut_reg[17]) );
  INVX16 U36 ( .A(n23), .Y(ALUOut_reg[18]) );
  INVX16 U37 ( .A(n22), .Y(ALUOut_reg[22]) );
  INVX16 U38 ( .A(n21), .Y(ALUOut_reg[23]) );
  INVX16 U39 ( .A(n20), .Y(ALUOut_reg[24]) );
  INVX16 U40 ( .A(n19), .Y(ALUOut_reg[28]) );
  INVX16 U41 ( .A(n18), .Y(ALUOut_reg[29]) );
  INVX16 U42 ( .A(n17), .Y(ALUOut_reg[30]) );
  INVX16 U43 ( .A(n16), .Y(ALUOut_reg[31]) );
  INVX16 U44 ( .A(n4), .Y(ALUOut_reg[7]) );
  INVX16 U45 ( .A(n3), .Y(ALUOut_reg[8]) );
  INVX16 U46 ( .A(n2), .Y(ALUOut_reg[9]) );
  INVX16 U47 ( .A(n1), .Y(ALUOut_reg[13]) );
  INVX16 U48 ( .A(n12), .Y(ALUOut_reg[14]) );
  INVX16 U49 ( .A(n11), .Y(ALUOut_reg[15]) );
  INVX16 U50 ( .A(n10), .Y(ALUOut_reg[19]) );
  INVX16 U51 ( .A(n9), .Y(ALUOut_reg[20]) );
  INVX16 U52 ( .A(n8), .Y(ALUOut_reg[21]) );
  INVX16 U53 ( .A(n7), .Y(ALUOut_reg[25]) );
  INVX16 U54 ( .A(n6), .Y(ALUOut_reg[26]) );
  INVX16 U55 ( .A(n5), .Y(ALUOut_reg[27]) );
  INVX16 U56 ( .A(n15), .Y(ALUOut_reg[10]) );
  INVX16 U57 ( .A(n14), .Y(ALUOut_reg[11]) );
  INVX16 U58 ( .A(n13), .Y(ALUOut_reg[12]) );
  BUFX16 U59 ( .A(n127), .Y(ALUOut_reg[3]) );
  BUFX16 U60 ( .A(n128), .Y(ALUOut_reg[2]) );
  INVX16 U61 ( .A(n117), .Y(M_reg[1]) );
  CLKBUFX3 U62 ( .A(stall_bothzero), .Y(n125) );
  CLKBUFX3 U63 ( .A(n120), .Y(n126) );
  CLKBUFX3 U64 ( .A(n120), .Y(n123) );
  CLKBUFX3 U65 ( .A(stall_bothzero), .Y(n122) );
  CLKBUFX3 U66 ( .A(stall_bothzero), .Y(n121) );
  CLKBUFX3 U67 ( .A(n120), .Y(n124) );
  CLKBUFX3 U68 ( .A(stall_bothzero), .Y(n120) );
  CLKBUFX3 U69 ( .A(stall_bothzero), .Y(n119) );
endmodule


module MEMWB ( clk, WB, Memout, ALUOut, RegRD, MEM_pcplus4, WBreg, Memreg, 
        ALUreg, RegRDreg, stall_bothzero, WB_pcplus4 );
  input [2:0] WB;
  input [31:0] Memout;
  input [31:0] ALUOut;
  input [4:0] RegRD;
  input [31:0] MEM_pcplus4;
  output [2:0] WBreg;
  output [31:0] Memreg;
  output [31:0] ALUreg;
  output [4:0] RegRDreg;
  output [31:0] WB_pcplus4;
  input clk, stall_bothzero;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  EDFFX1 \WB_pcplus4_reg[31]  ( .D(MEM_pcplus4[31]), .E(n1), .CK(clk), .Q(
        WB_pcplus4[31]) );
  EDFFX1 \WB_pcplus4_reg[30]  ( .D(MEM_pcplus4[30]), .E(n1), .CK(clk), .Q(
        WB_pcplus4[30]) );
  EDFFX1 \WB_pcplus4_reg[29]  ( .D(MEM_pcplus4[29]), .E(n1), .CK(clk), .Q(
        WB_pcplus4[29]) );
  EDFFX1 \WB_pcplus4_reg[28]  ( .D(MEM_pcplus4[28]), .E(n1), .CK(clk), .Q(
        WB_pcplus4[28]) );
  EDFFX1 \WB_pcplus4_reg[27]  ( .D(MEM_pcplus4[27]), .E(n1), .CK(clk), .Q(
        WB_pcplus4[27]) );
  EDFFX1 \WB_pcplus4_reg[26]  ( .D(MEM_pcplus4[26]), .E(n1), .CK(clk), .Q(
        WB_pcplus4[26]) );
  EDFFX1 \WB_pcplus4_reg[25]  ( .D(MEM_pcplus4[25]), .E(n2), .CK(clk), .Q(
        WB_pcplus4[25]) );
  EDFFX1 \WB_pcplus4_reg[24]  ( .D(MEM_pcplus4[24]), .E(n2), .CK(clk), .Q(
        WB_pcplus4[24]) );
  EDFFX1 \WB_pcplus4_reg[23]  ( .D(MEM_pcplus4[23]), .E(n2), .CK(clk), .Q(
        WB_pcplus4[23]) );
  EDFFX1 \WB_pcplus4_reg[22]  ( .D(MEM_pcplus4[22]), .E(n2), .CK(clk), .Q(
        WB_pcplus4[22]) );
  EDFFX1 \WB_pcplus4_reg[21]  ( .D(MEM_pcplus4[21]), .E(n2), .CK(clk), .Q(
        WB_pcplus4[21]) );
  EDFFX1 \WB_pcplus4_reg[20]  ( .D(MEM_pcplus4[20]), .E(n2), .CK(clk), .Q(
        WB_pcplus4[20]) );
  EDFFX1 \WB_pcplus4_reg[19]  ( .D(MEM_pcplus4[19]), .E(n2), .CK(clk), .Q(
        WB_pcplus4[19]) );
  EDFFX1 \WB_pcplus4_reg[18]  ( .D(MEM_pcplus4[18]), .E(n3), .CK(clk), .Q(
        WB_pcplus4[18]) );
  EDFFX1 \WB_pcplus4_reg[17]  ( .D(MEM_pcplus4[17]), .E(n3), .CK(clk), .Q(
        WB_pcplus4[17]) );
  EDFFX1 \WB_pcplus4_reg[16]  ( .D(MEM_pcplus4[16]), .E(n3), .CK(clk), .Q(
        WB_pcplus4[16]) );
  EDFFX1 \WB_pcplus4_reg[15]  ( .D(MEM_pcplus4[15]), .E(n3), .CK(clk), .Q(
        WB_pcplus4[15]) );
  EDFFX1 \WB_pcplus4_reg[14]  ( .D(MEM_pcplus4[14]), .E(n3), .CK(clk), .Q(
        WB_pcplus4[14]) );
  EDFFX1 \WB_pcplus4_reg[13]  ( .D(MEM_pcplus4[13]), .E(n3), .CK(clk), .Q(
        WB_pcplus4[13]) );
  EDFFX1 \WB_pcplus4_reg[12]  ( .D(MEM_pcplus4[12]), .E(n3), .CK(clk), .Q(
        WB_pcplus4[12]) );
  EDFFX1 \WB_pcplus4_reg[11]  ( .D(MEM_pcplus4[11]), .E(n4), .CK(clk), .Q(
        WB_pcplus4[11]) );
  EDFFX1 \WB_pcplus4_reg[10]  ( .D(MEM_pcplus4[10]), .E(n4), .CK(clk), .Q(
        WB_pcplus4[10]) );
  EDFFX1 \WB_pcplus4_reg[9]  ( .D(MEM_pcplus4[9]), .E(n4), .CK(clk), .Q(
        WB_pcplus4[9]) );
  EDFFX1 \WB_pcplus4_reg[8]  ( .D(MEM_pcplus4[8]), .E(n4), .CK(clk), .Q(
        WB_pcplus4[8]) );
  EDFFX1 \WB_pcplus4_reg[7]  ( .D(MEM_pcplus4[7]), .E(n4), .CK(clk), .Q(
        WB_pcplus4[7]) );
  EDFFX1 \WB_pcplus4_reg[6]  ( .D(MEM_pcplus4[6]), .E(n5), .CK(clk), .Q(
        WB_pcplus4[6]) );
  EDFFX1 \WB_pcplus4_reg[5]  ( .D(MEM_pcplus4[5]), .E(n5), .CK(clk), .Q(
        WB_pcplus4[5]) );
  EDFFX1 \WB_pcplus4_reg[4]  ( .D(MEM_pcplus4[4]), .E(n5), .CK(clk), .Q(
        WB_pcplus4[4]) );
  EDFFX1 \WB_pcplus4_reg[3]  ( .D(MEM_pcplus4[3]), .E(n5), .CK(clk), .Q(
        WB_pcplus4[3]) );
  EDFFX1 \WB_pcplus4_reg[2]  ( .D(MEM_pcplus4[2]), .E(n5), .CK(clk), .Q(
        WB_pcplus4[2]) );
  EDFFX1 \WB_pcplus4_reg[1]  ( .D(MEM_pcplus4[1]), .E(n8), .CK(clk), .Q(
        WB_pcplus4[1]) );
  EDFFX1 \WB_pcplus4_reg[0]  ( .D(MEM_pcplus4[0]), .E(n8), .CK(clk), .Q(
        WB_pcplus4[0]) );
  EDFFX1 \ALUreg_reg[31]  ( .D(ALUOut[31]), .E(n6), .CK(clk), .Q(ALUreg[31])
         );
  EDFFX1 \ALUreg_reg[30]  ( .D(ALUOut[30]), .E(n6), .CK(clk), .Q(ALUreg[30])
         );
  EDFFX1 \ALUreg_reg[29]  ( .D(ALUOut[29]), .E(n6), .CK(clk), .Q(ALUreg[29])
         );
  EDFFX1 \ALUreg_reg[28]  ( .D(ALUOut[28]), .E(n6), .CK(clk), .Q(ALUreg[28])
         );
  EDFFX1 \ALUreg_reg[27]  ( .D(ALUOut[27]), .E(n6), .CK(clk), .Q(ALUreg[27])
         );
  EDFFX1 \ALUreg_reg[26]  ( .D(ALUOut[26]), .E(n6), .CK(clk), .Q(ALUreg[26])
         );
  EDFFX1 \ALUreg_reg[25]  ( .D(ALUOut[25]), .E(n6), .CK(clk), .Q(ALUreg[25])
         );
  EDFFX1 \ALUreg_reg[24]  ( .D(ALUOut[24]), .E(n6), .CK(clk), .Q(ALUreg[24])
         );
  EDFFX1 \ALUreg_reg[23]  ( .D(ALUOut[23]), .E(n6), .CK(clk), .Q(ALUreg[23])
         );
  EDFFX1 \ALUreg_reg[22]  ( .D(ALUOut[22]), .E(n7), .CK(clk), .Q(ALUreg[22])
         );
  EDFFX1 \ALUreg_reg[21]  ( .D(ALUOut[21]), .E(n7), .CK(clk), .Q(ALUreg[21])
         );
  EDFFX1 \ALUreg_reg[20]  ( .D(ALUOut[20]), .E(n7), .CK(clk), .Q(ALUreg[20])
         );
  EDFFX1 \ALUreg_reg[19]  ( .D(ALUOut[19]), .E(n7), .CK(clk), .Q(ALUreg[19])
         );
  EDFFX1 \ALUreg_reg[18]  ( .D(ALUOut[18]), .E(n7), .CK(clk), .Q(ALUreg[18])
         );
  EDFFX1 \ALUreg_reg[17]  ( .D(ALUOut[17]), .E(n7), .CK(clk), .Q(ALUreg[17])
         );
  EDFFX1 \ALUreg_reg[16]  ( .D(ALUOut[16]), .E(n7), .CK(clk), .Q(ALUreg[16])
         );
  EDFFX1 \ALUreg_reg[15]  ( .D(ALUOut[15]), .E(n7), .CK(clk), .Q(ALUreg[15])
         );
  EDFFX1 \ALUreg_reg[14]  ( .D(ALUOut[14]), .E(n7), .CK(clk), .Q(ALUreg[14])
         );
  EDFFX1 \ALUreg_reg[13]  ( .D(ALUOut[13]), .E(n7), .CK(clk), .Q(ALUreg[13])
         );
  EDFFX1 \ALUreg_reg[12]  ( .D(ALUOut[12]), .E(n7), .CK(clk), .Q(ALUreg[12])
         );
  EDFFX1 \ALUreg_reg[11]  ( .D(ALUOut[11]), .E(n7), .CK(clk), .Q(ALUreg[11])
         );
  EDFFX1 \ALUreg_reg[10]  ( .D(ALUOut[10]), .E(n7), .CK(clk), .Q(ALUreg[10])
         );
  EDFFX1 \ALUreg_reg[9]  ( .D(ALUOut[9]), .E(n8), .CK(clk), .Q(ALUreg[9]) );
  EDFFX1 \ALUreg_reg[8]  ( .D(ALUOut[8]), .E(n8), .CK(clk), .Q(ALUreg[8]) );
  EDFFX1 \ALUreg_reg[7]  ( .D(ALUOut[7]), .E(n8), .CK(clk), .Q(ALUreg[7]) );
  EDFFX1 \ALUreg_reg[6]  ( .D(ALUOut[6]), .E(n8), .CK(clk), .Q(ALUreg[6]) );
  EDFFX1 \ALUreg_reg[5]  ( .D(ALUOut[5]), .E(n8), .CK(clk), .Q(ALUreg[5]) );
  EDFFX1 \ALUreg_reg[4]  ( .D(ALUOut[4]), .E(n8), .CK(clk), .Q(ALUreg[4]) );
  EDFFX1 \ALUreg_reg[3]  ( .D(ALUOut[3]), .E(n8), .CK(clk), .Q(ALUreg[3]) );
  EDFFX1 \ALUreg_reg[2]  ( .D(ALUOut[2]), .E(n8), .CK(clk), .Q(ALUreg[2]) );
  EDFFX1 \ALUreg_reg[1]  ( .D(ALUOut[1]), .E(n8), .CK(clk), .Q(ALUreg[1]) );
  EDFFX1 \ALUreg_reg[0]  ( .D(ALUOut[0]), .E(n8), .CK(clk), .Q(ALUreg[0]) );
  EDFFX1 \Memreg_reg[31]  ( .D(Memout[31]), .E(n1), .CK(clk), .Q(Memreg[31])
         );
  EDFFX1 \Memreg_reg[30]  ( .D(Memout[30]), .E(n1), .CK(clk), .Q(Memreg[30])
         );
  EDFFX1 \Memreg_reg[29]  ( .D(Memout[29]), .E(n1), .CK(clk), .Q(Memreg[29])
         );
  EDFFX1 \Memreg_reg[28]  ( .D(Memout[28]), .E(n1), .CK(clk), .Q(Memreg[28])
         );
  EDFFX1 \Memreg_reg[27]  ( .D(Memout[27]), .E(n1), .CK(clk), .Q(Memreg[27])
         );
  EDFFX1 \Memreg_reg[26]  ( .D(Memout[26]), .E(n1), .CK(clk), .Q(Memreg[26])
         );
  EDFFX1 \Memreg_reg[25]  ( .D(Memout[25]), .E(n1), .CK(clk), .Q(Memreg[25])
         );
  EDFFX1 \Memreg_reg[24]  ( .D(Memout[24]), .E(n2), .CK(clk), .Q(Memreg[24])
         );
  EDFFX1 \Memreg_reg[23]  ( .D(Memout[23]), .E(n2), .CK(clk), .Q(Memreg[23])
         );
  EDFFX1 \Memreg_reg[22]  ( .D(Memout[22]), .E(n2), .CK(clk), .Q(Memreg[22])
         );
  EDFFX1 \Memreg_reg[21]  ( .D(Memout[21]), .E(n2), .CK(clk), .Q(Memreg[21])
         );
  EDFFX1 \Memreg_reg[20]  ( .D(Memout[20]), .E(n2), .CK(clk), .Q(Memreg[20])
         );
  EDFFX1 \Memreg_reg[19]  ( .D(Memout[19]), .E(n2), .CK(clk), .Q(Memreg[19])
         );
  EDFFX1 \Memreg_reg[18]  ( .D(Memout[18]), .E(n8), .CK(clk), .Q(Memreg[18])
         );
  EDFFX1 \Memreg_reg[17]  ( .D(Memout[17]), .E(n3), .CK(clk), .Q(Memreg[17])
         );
  EDFFX1 \Memreg_reg[16]  ( .D(Memout[16]), .E(n3), .CK(clk), .Q(Memreg[16])
         );
  EDFFX1 \Memreg_reg[15]  ( .D(Memout[15]), .E(n3), .CK(clk), .Q(Memreg[15])
         );
  EDFFX1 \Memreg_reg[14]  ( .D(Memout[14]), .E(n3), .CK(clk), .Q(Memreg[14])
         );
  EDFFX1 \Memreg_reg[13]  ( .D(Memout[13]), .E(n3), .CK(clk), .Q(Memreg[13])
         );
  EDFFX1 \Memreg_reg[12]  ( .D(Memout[12]), .E(n3), .CK(clk), .Q(Memreg[12])
         );
  EDFFX1 \Memreg_reg[11]  ( .D(Memout[11]), .E(n4), .CK(clk), .Q(Memreg[11])
         );
  EDFFX1 \Memreg_reg[10]  ( .D(Memout[10]), .E(n4), .CK(clk), .Q(Memreg[10])
         );
  EDFFX1 \Memreg_reg[9]  ( .D(Memout[9]), .E(n4), .CK(clk), .Q(Memreg[9]) );
  EDFFX1 \Memreg_reg[8]  ( .D(Memout[8]), .E(n4), .CK(clk), .Q(Memreg[8]) );
  EDFFX1 \Memreg_reg[7]  ( .D(Memout[7]), .E(n4), .CK(clk), .Q(Memreg[7]) );
  EDFFX1 \Memreg_reg[6]  ( .D(Memout[6]), .E(n4), .CK(clk), .Q(Memreg[6]) );
  EDFFX1 \Memreg_reg[5]  ( .D(Memout[5]), .E(n4), .CK(clk), .Q(Memreg[5]) );
  EDFFX1 \Memreg_reg[4]  ( .D(Memout[4]), .E(n6), .CK(clk), .Q(Memreg[4]) );
  EDFFX1 \Memreg_reg[3]  ( .D(Memout[3]), .E(n6), .CK(clk), .Q(Memreg[3]) );
  EDFFX1 \Memreg_reg[2]  ( .D(Memout[2]), .E(n4), .CK(clk), .Q(Memreg[2]) );
  EDFFX1 \Memreg_reg[1]  ( .D(Memout[1]), .E(n5), .CK(clk), .Q(Memreg[1]) );
  EDFFX1 \Memreg_reg[0]  ( .D(Memout[0]), .E(n5), .CK(clk), .Q(Memreg[0]) );
  EDFFX1 \WBreg_reg[2]  ( .D(WB[2]), .E(n6), .CK(clk), .Q(WBreg[2]) );
  EDFFX1 \WBreg_reg[1]  ( .D(WB[1]), .E(n5), .CK(clk), .Q(WBreg[1]) );
  EDFFX1 \WBreg_reg[0]  ( .D(WB[0]), .E(n6), .CK(clk), .Q(WBreg[0]) );
  EDFFX1 \RegRDreg_reg[3]  ( .D(RegRD[3]), .E(n5), .CK(clk), .Q(RegRDreg[3])
         );
  EDFFX2 \RegRDreg_reg[4]  ( .D(RegRD[4]), .E(n5), .CK(clk), .Q(RegRDreg[4])
         );
  EDFFX2 \RegRDreg_reg[1]  ( .D(RegRD[1]), .E(n5), .CK(clk), .Q(RegRDreg[1])
         );
  EDFFX2 \RegRDreg_reg[0]  ( .D(RegRD[0]), .E(n5), .CK(clk), .Q(RegRDreg[0])
         );
  EDFFX2 \RegRDreg_reg[2]  ( .D(RegRD[2]), .E(n5), .CK(clk), .Q(RegRDreg[2])
         );
  CLKBUFX3 U2 ( .A(stall_bothzero), .Y(n7) );
  CLKBUFX3 U3 ( .A(stall_bothzero), .Y(n6) );
  CLKBUFX3 U4 ( .A(n3), .Y(n8) );
  CLKBUFX3 U5 ( .A(stall_bothzero), .Y(n4) );
  CLKBUFX3 U6 ( .A(stall_bothzero), .Y(n3) );
  CLKBUFX3 U7 ( .A(stall_bothzero), .Y(n2) );
  CLKBUFX3 U8 ( .A(stall_bothzero), .Y(n1) );
  CLKBUFX3 U9 ( .A(stall_bothzero), .Y(n5) );
endmodule


module MIPS_Pipeline_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  XOR3XL U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  AND2X2 U1 ( .A(B[2]), .B(A[2]), .Y(n1) );
  XOR2X1 U2 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  BUFX2 U3 ( .A(A[0]), .Y(SUM[0]) );
  BUFX2 U4 ( .A(A[1]), .Y(SUM[1]) );
endmodule


module MIPS_Pipeline_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  CLKINVX1 U1 ( .A(B[1]), .Y(n2) );
  CLKINVX1 U2 ( .A(A[1]), .Y(n1) );
  NOR4X1 U3 ( .A(n3), .B(n4), .C(n5), .D(n6), .Y(EQ) );
  NAND4X1 U4 ( .A(n7), .B(n8), .C(n9), .D(n10), .Y(n6) );
  XNOR2X1 U5 ( .A(B[11]), .B(A[11]), .Y(n10) );
  XNOR2X1 U6 ( .A(B[12]), .B(A[12]), .Y(n9) );
  XNOR2X1 U7 ( .A(B[13]), .B(A[13]), .Y(n8) );
  XNOR2X1 U8 ( .A(B[14]), .B(A[14]), .Y(n7) );
  NAND4X1 U9 ( .A(n11), .B(n12), .C(n13), .D(n14), .Y(n5) );
  XNOR2X1 U10 ( .A(B[7]), .B(A[7]), .Y(n14) );
  XNOR2X1 U11 ( .A(B[8]), .B(A[8]), .Y(n13) );
  XNOR2X1 U12 ( .A(B[9]), .B(A[9]), .Y(n12) );
  XNOR2X1 U13 ( .A(B[10]), .B(A[10]), .Y(n11) );
  NAND4X1 U14 ( .A(n15), .B(n16), .C(n17), .D(n18), .Y(n4) );
  NOR4X1 U15 ( .A(n19), .B(n20), .C(n21), .D(n22), .Y(n18) );
  XOR2X1 U16 ( .A(B[6]), .B(A[6]), .Y(n22) );
  XOR2X1 U17 ( .A(B[5]), .B(A[5]), .Y(n21) );
  XOR2X1 U18 ( .A(B[4]), .B(A[4]), .Y(n20) );
  XOR2X1 U19 ( .A(B[3]), .B(A[3]), .Y(n19) );
  NOR2X1 U20 ( .A(n23), .B(n24), .Y(n17) );
  XOR2X1 U21 ( .A(B[2]), .B(A[2]), .Y(n24) );
  XOR2X1 U22 ( .A(B[31]), .B(A[31]), .Y(n23) );
  OAI22XL U23 ( .A0(n25), .A1(n1), .B0(B[1]), .B1(n25), .Y(n16) );
  NOR2BX1 U24 ( .AN(B[0]), .B(A[0]), .Y(n25) );
  OAI22XL U25 ( .A0(A[1]), .A1(n26), .B0(n26), .B1(n2), .Y(n15) );
  NOR2BX1 U26 ( .AN(A[0]), .B(B[0]), .Y(n26) );
  NAND4X1 U27 ( .A(n27), .B(n28), .C(n29), .D(n30), .Y(n3) );
  NOR4X1 U28 ( .A(n31), .B(n32), .C(n33), .D(n34), .Y(n30) );
  XOR2X1 U29 ( .A(B[18]), .B(A[18]), .Y(n34) );
  XOR2X1 U30 ( .A(B[17]), .B(A[17]), .Y(n33) );
  XOR2X1 U31 ( .A(B[16]), .B(A[16]), .Y(n32) );
  XOR2X1 U32 ( .A(B[15]), .B(A[15]), .Y(n31) );
  NOR4X1 U33 ( .A(n35), .B(n36), .C(n37), .D(n38), .Y(n29) );
  XOR2X1 U34 ( .A(B[22]), .B(A[22]), .Y(n38) );
  XOR2X1 U35 ( .A(B[21]), .B(A[21]), .Y(n37) );
  XOR2X1 U36 ( .A(B[20]), .B(A[20]), .Y(n36) );
  XOR2X1 U37 ( .A(B[19]), .B(A[19]), .Y(n35) );
  NOR4X1 U38 ( .A(n39), .B(n40), .C(n41), .D(n42), .Y(n28) );
  XOR2X1 U39 ( .A(B[26]), .B(A[26]), .Y(n42) );
  XOR2X1 U40 ( .A(B[25]), .B(A[25]), .Y(n41) );
  XOR2X1 U41 ( .A(B[24]), .B(A[24]), .Y(n40) );
  XOR2X1 U42 ( .A(B[23]), .B(A[23]), .Y(n39) );
  NOR4X1 U43 ( .A(n43), .B(n44), .C(n45), .D(n46), .Y(n27) );
  XOR2X1 U44 ( .A(B[30]), .B(A[30]), .Y(n46) );
  XOR2X1 U45 ( .A(B[29]), .B(A[29]), .Y(n45) );
  XOR2X1 U46 ( .A(B[28]), .B(A[28]), .Y(n44) );
  XOR2X1 U47 ( .A(B[27]), .B(A[27]), .Y(n43) );
endmodule


module MIPS_Pipeline_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n30;

  XOR2X1 U1 ( .A(A[3]), .B(A[2]), .Y(SUM[3]) );
  XOR2X1 U2 ( .A(A[7]), .B(n1), .Y(SUM[7]) );
  XOR2X1 U3 ( .A(A[4]), .B(n2), .Y(SUM[4]) );
  XOR2X1 U4 ( .A(A[5]), .B(n3), .Y(SUM[5]) );
  XOR2X1 U5 ( .A(A[6]), .B(n4), .Y(SUM[6]) );
  XOR2X1 U6 ( .A(A[8]), .B(n5), .Y(SUM[8]) );
  XOR2X1 U7 ( .A(A[9]), .B(n6), .Y(SUM[9]) );
  XOR2X1 U8 ( .A(A[10]), .B(n7), .Y(SUM[10]) );
  XOR2X1 U9 ( .A(A[11]), .B(n17), .Y(SUM[11]) );
  XOR2X1 U10 ( .A(A[12]), .B(n18), .Y(SUM[12]) );
  XOR2X1 U11 ( .A(A[13]), .B(n19), .Y(SUM[13]) );
  XOR2X1 U12 ( .A(A[14]), .B(n8), .Y(SUM[14]) );
  XOR2X1 U13 ( .A(A[15]), .B(n9), .Y(SUM[15]) );
  XOR2X1 U14 ( .A(A[16]), .B(n10), .Y(SUM[16]) );
  XOR2X1 U15 ( .A(A[17]), .B(n20), .Y(SUM[17]) );
  XOR2X1 U16 ( .A(A[18]), .B(n21), .Y(SUM[18]) );
  XOR2X1 U17 ( .A(A[19]), .B(n22), .Y(SUM[19]) );
  XOR2X1 U18 ( .A(A[20]), .B(n11), .Y(SUM[20]) );
  XOR2X1 U19 ( .A(A[21]), .B(n12), .Y(SUM[21]) );
  XOR2X1 U20 ( .A(A[22]), .B(n13), .Y(SUM[22]) );
  XOR2X1 U21 ( .A(A[23]), .B(n23), .Y(SUM[23]) );
  XOR2X1 U22 ( .A(A[24]), .B(n24), .Y(SUM[24]) );
  XOR2X1 U23 ( .A(A[25]), .B(n25), .Y(SUM[25]) );
  XOR2X1 U24 ( .A(A[26]), .B(n14), .Y(SUM[26]) );
  XOR2X1 U25 ( .A(A[27]), .B(n15), .Y(SUM[27]) );
  XOR2X1 U26 ( .A(A[28]), .B(n16), .Y(SUM[28]) );
  XOR2X1 U27 ( .A(A[29]), .B(n26), .Y(SUM[29]) );
  XOR2X1 U28 ( .A(A[30]), .B(n27), .Y(SUM[30]) );
  XNOR2X1 U29 ( .A(A[31]), .B(n30), .Y(SUM[31]) );
  NAND2X1 U30 ( .A(A[30]), .B(n27), .Y(n30) );
  CLKINVX1 U31 ( .A(A[2]), .Y(SUM[2]) );
  AND2X2 U32 ( .A(A[6]), .B(n4), .Y(n1) );
  AND2X2 U33 ( .A(A[3]), .B(A[2]), .Y(n2) );
  AND2X2 U34 ( .A(A[4]), .B(n2), .Y(n3) );
  AND2X2 U35 ( .A(A[5]), .B(n3), .Y(n4) );
  AND2X2 U36 ( .A(A[7]), .B(n1), .Y(n5) );
  AND2X2 U37 ( .A(A[8]), .B(n5), .Y(n6) );
  AND2X2 U38 ( .A(A[9]), .B(n6), .Y(n7) );
  AND2X2 U39 ( .A(A[13]), .B(n19), .Y(n8) );
  AND2X2 U40 ( .A(A[14]), .B(n8), .Y(n9) );
  AND2X2 U41 ( .A(A[15]), .B(n9), .Y(n10) );
  AND2X2 U42 ( .A(A[19]), .B(n22), .Y(n11) );
  AND2X2 U43 ( .A(A[20]), .B(n11), .Y(n12) );
  AND2X2 U44 ( .A(A[21]), .B(n12), .Y(n13) );
  AND2X2 U45 ( .A(A[25]), .B(n25), .Y(n14) );
  AND2X2 U46 ( .A(A[26]), .B(n14), .Y(n15) );
  AND2X2 U47 ( .A(A[27]), .B(n15), .Y(n16) );
  AND2X2 U48 ( .A(A[10]), .B(n7), .Y(n17) );
  AND2X2 U49 ( .A(A[11]), .B(n17), .Y(n18) );
  AND2X2 U50 ( .A(A[12]), .B(n18), .Y(n19) );
  AND2X2 U51 ( .A(A[16]), .B(n10), .Y(n20) );
  AND2X2 U52 ( .A(A[17]), .B(n20), .Y(n21) );
  AND2X2 U53 ( .A(A[18]), .B(n21), .Y(n22) );
  AND2X2 U54 ( .A(A[22]), .B(n13), .Y(n23) );
  AND2X2 U55 ( .A(A[23]), .B(n23), .Y(n24) );
  AND2X2 U56 ( .A(A[24]), .B(n24), .Y(n25) );
  AND2X2 U57 ( .A(A[28]), .B(n16), .Y(n26) );
  AND2X2 U58 ( .A(A[29]), .B(n26), .Y(n27) );
  BUFX2 U59 ( .A(A[0]), .Y(SUM[0]) );
  BUFX2 U60 ( .A(A[1]), .Y(SUM[1]) );
endmodule


module MIPS_Pipeline ( clk, rst_n, ICACHE_ren, ICACHE_wen, ICACHE_addr, 
        ICACHE_wdata, ICACHE_stall, ICACHE_rdata, DCACHE_ren, DCACHE_wen, 
        DCACHE_addr, DCACHE_wdata, DCACHE_stall, DCACHE_rdata );
  output [29:0] ICACHE_addr;
  output [31:0] ICACHE_wdata;
  input [31:0] ICACHE_rdata;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input [31:0] DCACHE_rdata;
  input clk, rst_n, ICACHE_stall, DCACHE_stall;
  output ICACHE_ren, ICACHE_wen, DCACHE_ren, DCACHE_wen;
  wire   N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, IFIDWrite, PCWrite,
         \MemtoReg[0] , \reg_file_next[0][31] , \reg_file_next[0][30] ,
         \reg_file_next[0][29] , \reg_file_next[0][28] ,
         \reg_file_next[0][27] , \reg_file_next[0][26] ,
         \reg_file_next[0][25] , \reg_file_next[0][24] ,
         \reg_file_next[0][23] , \reg_file_next[0][22] ,
         \reg_file_next[0][21] , \reg_file_next[0][20] ,
         \reg_file_next[0][19] , \reg_file_next[0][18] ,
         \reg_file_next[0][17] , \reg_file_next[0][16] ,
         \reg_file_next[0][15] , \reg_file_next[0][14] ,
         \reg_file_next[0][13] , \reg_file_next[0][12] ,
         \reg_file_next[0][11] , \reg_file_next[0][10] , \reg_file_next[0][9] ,
         \reg_file_next[0][8] , \reg_file_next[0][7] , \reg_file_next[0][6] ,
         \reg_file_next[0][5] , \reg_file_next[0][4] , \reg_file_next[0][3] ,
         \reg_file_next[0][2] , \reg_file_next[0][1] , \reg_file_next[0][0] ,
         \reg_file_next[1][31] , \reg_file_next[1][30] ,
         \reg_file_next[1][29] , \reg_file_next[1][28] ,
         \reg_file_next[1][27] , \reg_file_next[1][26] ,
         \reg_file_next[1][25] , \reg_file_next[1][24] ,
         \reg_file_next[1][23] , \reg_file_next[1][22] ,
         \reg_file_next[1][21] , \reg_file_next[1][20] ,
         \reg_file_next[1][19] , \reg_file_next[1][18] ,
         \reg_file_next[1][17] , \reg_file_next[1][16] ,
         \reg_file_next[1][15] , \reg_file_next[1][14] ,
         \reg_file_next[1][13] , \reg_file_next[1][12] ,
         \reg_file_next[1][11] , \reg_file_next[1][10] , \reg_file_next[1][9] ,
         \reg_file_next[1][8] , \reg_file_next[1][7] , \reg_file_next[1][6] ,
         \reg_file_next[1][5] , \reg_file_next[1][4] , \reg_file_next[1][3] ,
         \reg_file_next[1][2] , \reg_file_next[1][1] , \reg_file_next[1][0] ,
         \reg_file_next[2][31] , \reg_file_next[2][30] ,
         \reg_file_next[2][29] , \reg_file_next[2][28] ,
         \reg_file_next[2][27] , \reg_file_next[2][26] ,
         \reg_file_next[2][25] , \reg_file_next[2][24] ,
         \reg_file_next[2][23] , \reg_file_next[2][22] ,
         \reg_file_next[2][21] , \reg_file_next[2][20] ,
         \reg_file_next[2][19] , \reg_file_next[2][18] ,
         \reg_file_next[2][17] , \reg_file_next[2][16] ,
         \reg_file_next[2][15] , \reg_file_next[2][14] ,
         \reg_file_next[2][13] , \reg_file_next[2][12] ,
         \reg_file_next[2][11] , \reg_file_next[2][10] , \reg_file_next[2][9] ,
         \reg_file_next[2][8] , \reg_file_next[2][7] , \reg_file_next[2][6] ,
         \reg_file_next[2][5] , \reg_file_next[2][4] , \reg_file_next[2][3] ,
         \reg_file_next[2][2] , \reg_file_next[2][1] , \reg_file_next[2][0] ,
         \reg_file_next[3][31] , \reg_file_next[3][30] ,
         \reg_file_next[3][29] , \reg_file_next[3][28] ,
         \reg_file_next[3][27] , \reg_file_next[3][26] ,
         \reg_file_next[3][25] , \reg_file_next[3][24] ,
         \reg_file_next[3][23] , \reg_file_next[3][22] ,
         \reg_file_next[3][21] , \reg_file_next[3][20] ,
         \reg_file_next[3][19] , \reg_file_next[3][18] ,
         \reg_file_next[3][17] , \reg_file_next[3][16] ,
         \reg_file_next[3][15] , \reg_file_next[3][14] ,
         \reg_file_next[3][13] , \reg_file_next[3][12] ,
         \reg_file_next[3][11] , \reg_file_next[3][10] , \reg_file_next[3][9] ,
         \reg_file_next[3][8] , \reg_file_next[3][7] , \reg_file_next[3][6] ,
         \reg_file_next[3][5] , \reg_file_next[3][4] , \reg_file_next[3][3] ,
         \reg_file_next[3][2] , \reg_file_next[3][1] , \reg_file_next[3][0] ,
         \reg_file_next[4][31] , \reg_file_next[4][30] ,
         \reg_file_next[4][29] , \reg_file_next[4][28] ,
         \reg_file_next[4][27] , \reg_file_next[4][26] ,
         \reg_file_next[4][25] , \reg_file_next[4][24] ,
         \reg_file_next[4][23] , \reg_file_next[4][22] ,
         \reg_file_next[4][21] , \reg_file_next[4][20] ,
         \reg_file_next[4][19] , \reg_file_next[4][18] ,
         \reg_file_next[4][17] , \reg_file_next[4][16] ,
         \reg_file_next[4][15] , \reg_file_next[4][14] ,
         \reg_file_next[4][13] , \reg_file_next[4][12] ,
         \reg_file_next[4][11] , \reg_file_next[4][10] , \reg_file_next[4][9] ,
         \reg_file_next[4][8] , \reg_file_next[4][7] , \reg_file_next[4][6] ,
         \reg_file_next[4][5] , \reg_file_next[4][4] , \reg_file_next[4][3] ,
         \reg_file_next[4][2] , \reg_file_next[4][1] , \reg_file_next[4][0] ,
         \reg_file_next[5][31] , \reg_file_next[5][30] ,
         \reg_file_next[5][29] , \reg_file_next[5][28] ,
         \reg_file_next[5][27] , \reg_file_next[5][26] ,
         \reg_file_next[5][25] , \reg_file_next[5][24] ,
         \reg_file_next[5][23] , \reg_file_next[5][22] ,
         \reg_file_next[5][21] , \reg_file_next[5][20] ,
         \reg_file_next[5][19] , \reg_file_next[5][18] ,
         \reg_file_next[5][17] , \reg_file_next[5][16] ,
         \reg_file_next[5][15] , \reg_file_next[5][14] ,
         \reg_file_next[5][13] , \reg_file_next[5][12] ,
         \reg_file_next[5][11] , \reg_file_next[5][10] , \reg_file_next[5][9] ,
         \reg_file_next[5][8] , \reg_file_next[5][7] , \reg_file_next[5][6] ,
         \reg_file_next[5][5] , \reg_file_next[5][4] , \reg_file_next[5][3] ,
         \reg_file_next[5][2] , \reg_file_next[5][1] , \reg_file_next[5][0] ,
         \reg_file_next[6][31] , \reg_file_next[6][30] ,
         \reg_file_next[6][29] , \reg_file_next[6][28] ,
         \reg_file_next[6][27] , \reg_file_next[6][26] ,
         \reg_file_next[6][25] , \reg_file_next[6][24] ,
         \reg_file_next[6][23] , \reg_file_next[6][22] ,
         \reg_file_next[6][21] , \reg_file_next[6][20] ,
         \reg_file_next[6][19] , \reg_file_next[6][18] ,
         \reg_file_next[6][17] , \reg_file_next[6][16] ,
         \reg_file_next[6][15] , \reg_file_next[6][14] ,
         \reg_file_next[6][13] , \reg_file_next[6][12] ,
         \reg_file_next[6][11] , \reg_file_next[6][10] , \reg_file_next[6][9] ,
         \reg_file_next[6][8] , \reg_file_next[6][7] , \reg_file_next[6][6] ,
         \reg_file_next[6][5] , \reg_file_next[6][4] , \reg_file_next[6][3] ,
         \reg_file_next[6][2] , \reg_file_next[6][1] , \reg_file_next[6][0] ,
         \reg_file_next[7][31] , \reg_file_next[7][30] ,
         \reg_file_next[7][29] , \reg_file_next[7][28] ,
         \reg_file_next[7][27] , \reg_file_next[7][26] ,
         \reg_file_next[7][25] , \reg_file_next[7][24] ,
         \reg_file_next[7][23] , \reg_file_next[7][22] ,
         \reg_file_next[7][21] , \reg_file_next[7][20] ,
         \reg_file_next[7][19] , \reg_file_next[7][18] ,
         \reg_file_next[7][17] , \reg_file_next[7][16] ,
         \reg_file_next[7][15] , \reg_file_next[7][14] ,
         \reg_file_next[7][13] , \reg_file_next[7][12] ,
         \reg_file_next[7][11] , \reg_file_next[7][10] , \reg_file_next[7][9] ,
         \reg_file_next[7][8] , \reg_file_next[7][7] , \reg_file_next[7][6] ,
         \reg_file_next[7][5] , \reg_file_next[7][4] , \reg_file_next[7][3] ,
         \reg_file_next[7][2] , \reg_file_next[7][1] , \reg_file_next[7][0] ,
         \reg_file_next[8][31] , \reg_file_next[8][30] ,
         \reg_file_next[8][29] , \reg_file_next[8][28] ,
         \reg_file_next[8][27] , \reg_file_next[8][26] ,
         \reg_file_next[8][25] , \reg_file_next[8][24] ,
         \reg_file_next[8][23] , \reg_file_next[8][22] ,
         \reg_file_next[8][21] , \reg_file_next[8][20] ,
         \reg_file_next[8][19] , \reg_file_next[8][18] ,
         \reg_file_next[8][17] , \reg_file_next[8][16] ,
         \reg_file_next[8][15] , \reg_file_next[8][14] ,
         \reg_file_next[8][13] , \reg_file_next[8][12] ,
         \reg_file_next[8][11] , \reg_file_next[8][10] , \reg_file_next[8][9] ,
         \reg_file_next[8][8] , \reg_file_next[8][7] , \reg_file_next[8][6] ,
         \reg_file_next[8][5] , \reg_file_next[8][4] , \reg_file_next[8][3] ,
         \reg_file_next[8][2] , \reg_file_next[8][1] , \reg_file_next[8][0] ,
         \reg_file_next[9][31] , \reg_file_next[9][30] ,
         \reg_file_next[9][29] , \reg_file_next[9][28] ,
         \reg_file_next[9][27] , \reg_file_next[9][26] ,
         \reg_file_next[9][25] , \reg_file_next[9][24] ,
         \reg_file_next[9][23] , \reg_file_next[9][22] ,
         \reg_file_next[9][21] , \reg_file_next[9][20] ,
         \reg_file_next[9][19] , \reg_file_next[9][18] ,
         \reg_file_next[9][17] , \reg_file_next[9][16] ,
         \reg_file_next[9][15] , \reg_file_next[9][14] ,
         \reg_file_next[9][13] , \reg_file_next[9][12] ,
         \reg_file_next[9][11] , \reg_file_next[9][10] , \reg_file_next[9][9] ,
         \reg_file_next[9][8] , \reg_file_next[9][7] , \reg_file_next[9][6] ,
         \reg_file_next[9][5] , \reg_file_next[9][4] , \reg_file_next[9][3] ,
         \reg_file_next[9][2] , \reg_file_next[9][1] , \reg_file_next[9][0] ,
         \reg_file_next[10][31] , \reg_file_next[10][30] ,
         \reg_file_next[10][29] , \reg_file_next[10][28] ,
         \reg_file_next[10][27] , \reg_file_next[10][26] ,
         \reg_file_next[10][25] , \reg_file_next[10][24] ,
         \reg_file_next[10][23] , \reg_file_next[10][22] ,
         \reg_file_next[10][21] , \reg_file_next[10][20] ,
         \reg_file_next[10][19] , \reg_file_next[10][18] ,
         \reg_file_next[10][17] , \reg_file_next[10][16] ,
         \reg_file_next[10][15] , \reg_file_next[10][14] ,
         \reg_file_next[10][13] , \reg_file_next[10][12] ,
         \reg_file_next[10][11] , \reg_file_next[10][10] ,
         \reg_file_next[10][9] , \reg_file_next[10][8] ,
         \reg_file_next[10][7] , \reg_file_next[10][6] ,
         \reg_file_next[10][5] , \reg_file_next[10][4] ,
         \reg_file_next[10][3] , \reg_file_next[10][2] ,
         \reg_file_next[10][1] , \reg_file_next[10][0] ,
         \reg_file_next[11][31] , \reg_file_next[11][30] ,
         \reg_file_next[11][29] , \reg_file_next[11][28] ,
         \reg_file_next[11][27] , \reg_file_next[11][26] ,
         \reg_file_next[11][25] , \reg_file_next[11][24] ,
         \reg_file_next[11][23] , \reg_file_next[11][22] ,
         \reg_file_next[11][21] , \reg_file_next[11][20] ,
         \reg_file_next[11][19] , \reg_file_next[11][18] ,
         \reg_file_next[11][17] , \reg_file_next[11][16] ,
         \reg_file_next[11][15] , \reg_file_next[11][14] ,
         \reg_file_next[11][13] , \reg_file_next[11][12] ,
         \reg_file_next[11][11] , \reg_file_next[11][10] ,
         \reg_file_next[11][9] , \reg_file_next[11][8] ,
         \reg_file_next[11][7] , \reg_file_next[11][6] ,
         \reg_file_next[11][5] , \reg_file_next[11][4] ,
         \reg_file_next[11][3] , \reg_file_next[11][2] ,
         \reg_file_next[11][1] , \reg_file_next[11][0] ,
         \reg_file_next[12][31] , \reg_file_next[12][30] ,
         \reg_file_next[12][29] , \reg_file_next[12][28] ,
         \reg_file_next[12][27] , \reg_file_next[12][26] ,
         \reg_file_next[12][25] , \reg_file_next[12][24] ,
         \reg_file_next[12][23] , \reg_file_next[12][22] ,
         \reg_file_next[12][21] , \reg_file_next[12][20] ,
         \reg_file_next[12][19] , \reg_file_next[12][18] ,
         \reg_file_next[12][17] , \reg_file_next[12][16] ,
         \reg_file_next[12][15] , \reg_file_next[12][14] ,
         \reg_file_next[12][13] , \reg_file_next[12][12] ,
         \reg_file_next[12][11] , \reg_file_next[12][10] ,
         \reg_file_next[12][9] , \reg_file_next[12][8] ,
         \reg_file_next[12][7] , \reg_file_next[12][6] ,
         \reg_file_next[12][5] , \reg_file_next[12][4] ,
         \reg_file_next[12][3] , \reg_file_next[12][2] ,
         \reg_file_next[12][1] , \reg_file_next[12][0] ,
         \reg_file_next[13][31] , \reg_file_next[13][30] ,
         \reg_file_next[13][29] , \reg_file_next[13][28] ,
         \reg_file_next[13][27] , \reg_file_next[13][26] ,
         \reg_file_next[13][25] , \reg_file_next[13][24] ,
         \reg_file_next[13][23] , \reg_file_next[13][22] ,
         \reg_file_next[13][21] , \reg_file_next[13][20] ,
         \reg_file_next[13][19] , \reg_file_next[13][18] ,
         \reg_file_next[13][17] , \reg_file_next[13][16] ,
         \reg_file_next[13][15] , \reg_file_next[13][14] ,
         \reg_file_next[13][13] , \reg_file_next[13][12] ,
         \reg_file_next[13][11] , \reg_file_next[13][10] ,
         \reg_file_next[13][9] , \reg_file_next[13][8] ,
         \reg_file_next[13][7] , \reg_file_next[13][6] ,
         \reg_file_next[13][5] , \reg_file_next[13][4] ,
         \reg_file_next[13][3] , \reg_file_next[13][2] ,
         \reg_file_next[13][1] , \reg_file_next[13][0] ,
         \reg_file_next[14][31] , \reg_file_next[14][30] ,
         \reg_file_next[14][29] , \reg_file_next[14][28] ,
         \reg_file_next[14][27] , \reg_file_next[14][26] ,
         \reg_file_next[14][25] , \reg_file_next[14][24] ,
         \reg_file_next[14][23] , \reg_file_next[14][22] ,
         \reg_file_next[14][21] , \reg_file_next[14][20] ,
         \reg_file_next[14][19] , \reg_file_next[14][18] ,
         \reg_file_next[14][17] , \reg_file_next[14][16] ,
         \reg_file_next[14][15] , \reg_file_next[14][14] ,
         \reg_file_next[14][13] , \reg_file_next[14][12] ,
         \reg_file_next[14][11] , \reg_file_next[14][10] ,
         \reg_file_next[14][9] , \reg_file_next[14][8] ,
         \reg_file_next[14][7] , \reg_file_next[14][6] ,
         \reg_file_next[14][5] , \reg_file_next[14][4] ,
         \reg_file_next[14][3] , \reg_file_next[14][2] ,
         \reg_file_next[14][1] , \reg_file_next[14][0] ,
         \reg_file_next[15][31] , \reg_file_next[15][30] ,
         \reg_file_next[15][29] , \reg_file_next[15][28] ,
         \reg_file_next[15][27] , \reg_file_next[15][26] ,
         \reg_file_next[15][25] , \reg_file_next[15][24] ,
         \reg_file_next[15][23] , \reg_file_next[15][22] ,
         \reg_file_next[15][21] , \reg_file_next[15][20] ,
         \reg_file_next[15][19] , \reg_file_next[15][18] ,
         \reg_file_next[15][17] , \reg_file_next[15][16] ,
         \reg_file_next[15][15] , \reg_file_next[15][14] ,
         \reg_file_next[15][13] , \reg_file_next[15][12] ,
         \reg_file_next[15][11] , \reg_file_next[15][10] ,
         \reg_file_next[15][9] , \reg_file_next[15][8] ,
         \reg_file_next[15][7] , \reg_file_next[15][6] ,
         \reg_file_next[15][5] , \reg_file_next[15][4] ,
         \reg_file_next[15][3] , \reg_file_next[15][2] ,
         \reg_file_next[15][1] , \reg_file_next[15][0] ,
         \reg_file_next[16][31] , \reg_file_next[16][30] ,
         \reg_file_next[16][29] , \reg_file_next[16][28] ,
         \reg_file_next[16][27] , \reg_file_next[16][26] ,
         \reg_file_next[16][25] , \reg_file_next[16][24] ,
         \reg_file_next[16][23] , \reg_file_next[16][22] ,
         \reg_file_next[16][21] , \reg_file_next[16][20] ,
         \reg_file_next[16][19] , \reg_file_next[16][18] ,
         \reg_file_next[16][17] , \reg_file_next[16][16] ,
         \reg_file_next[16][15] , \reg_file_next[16][14] ,
         \reg_file_next[16][13] , \reg_file_next[16][12] ,
         \reg_file_next[16][11] , \reg_file_next[16][10] ,
         \reg_file_next[16][9] , \reg_file_next[16][8] ,
         \reg_file_next[16][7] , \reg_file_next[16][6] ,
         \reg_file_next[16][5] , \reg_file_next[16][4] ,
         \reg_file_next[16][3] , \reg_file_next[16][2] ,
         \reg_file_next[16][1] , \reg_file_next[16][0] ,
         \reg_file_next[17][31] , \reg_file_next[17][30] ,
         \reg_file_next[17][29] , \reg_file_next[17][28] ,
         \reg_file_next[17][27] , \reg_file_next[17][26] ,
         \reg_file_next[17][25] , \reg_file_next[17][24] ,
         \reg_file_next[17][23] , \reg_file_next[17][22] ,
         \reg_file_next[17][21] , \reg_file_next[17][20] ,
         \reg_file_next[17][19] , \reg_file_next[17][18] ,
         \reg_file_next[17][17] , \reg_file_next[17][16] ,
         \reg_file_next[17][15] , \reg_file_next[17][14] ,
         \reg_file_next[17][13] , \reg_file_next[17][12] ,
         \reg_file_next[17][11] , \reg_file_next[17][10] ,
         \reg_file_next[17][9] , \reg_file_next[17][8] ,
         \reg_file_next[17][7] , \reg_file_next[17][6] ,
         \reg_file_next[17][5] , \reg_file_next[17][4] ,
         \reg_file_next[17][3] , \reg_file_next[17][2] ,
         \reg_file_next[17][1] , \reg_file_next[17][0] ,
         \reg_file_next[18][31] , \reg_file_next[18][30] ,
         \reg_file_next[18][29] , \reg_file_next[18][28] ,
         \reg_file_next[18][27] , \reg_file_next[18][26] ,
         \reg_file_next[18][25] , \reg_file_next[18][24] ,
         \reg_file_next[18][23] , \reg_file_next[18][22] ,
         \reg_file_next[18][21] , \reg_file_next[18][20] ,
         \reg_file_next[18][19] , \reg_file_next[18][18] ,
         \reg_file_next[18][17] , \reg_file_next[18][16] ,
         \reg_file_next[18][15] , \reg_file_next[18][14] ,
         \reg_file_next[18][13] , \reg_file_next[18][12] ,
         \reg_file_next[18][11] , \reg_file_next[18][10] ,
         \reg_file_next[18][9] , \reg_file_next[18][8] ,
         \reg_file_next[18][7] , \reg_file_next[18][6] ,
         \reg_file_next[18][5] , \reg_file_next[18][4] ,
         \reg_file_next[18][3] , \reg_file_next[18][2] ,
         \reg_file_next[18][1] , \reg_file_next[18][0] ,
         \reg_file_next[19][31] , \reg_file_next[19][30] ,
         \reg_file_next[19][29] , \reg_file_next[19][28] ,
         \reg_file_next[19][27] , \reg_file_next[19][26] ,
         \reg_file_next[19][25] , \reg_file_next[19][24] ,
         \reg_file_next[19][23] , \reg_file_next[19][22] ,
         \reg_file_next[19][21] , \reg_file_next[19][20] ,
         \reg_file_next[19][19] , \reg_file_next[19][18] ,
         \reg_file_next[19][17] , \reg_file_next[19][16] ,
         \reg_file_next[19][15] , \reg_file_next[19][14] ,
         \reg_file_next[19][13] , \reg_file_next[19][12] ,
         \reg_file_next[19][11] , \reg_file_next[19][10] ,
         \reg_file_next[19][9] , \reg_file_next[19][8] ,
         \reg_file_next[19][7] , \reg_file_next[19][6] ,
         \reg_file_next[19][5] , \reg_file_next[19][4] ,
         \reg_file_next[19][3] , \reg_file_next[19][2] ,
         \reg_file_next[19][1] , \reg_file_next[19][0] ,
         \reg_file_next[20][31] , \reg_file_next[20][30] ,
         \reg_file_next[20][29] , \reg_file_next[20][28] ,
         \reg_file_next[20][27] , \reg_file_next[20][26] ,
         \reg_file_next[20][25] , \reg_file_next[20][24] ,
         \reg_file_next[20][23] , \reg_file_next[20][22] ,
         \reg_file_next[20][21] , \reg_file_next[20][20] ,
         \reg_file_next[20][19] , \reg_file_next[20][18] ,
         \reg_file_next[20][17] , \reg_file_next[20][16] ,
         \reg_file_next[20][15] , \reg_file_next[20][14] ,
         \reg_file_next[20][13] , \reg_file_next[20][12] ,
         \reg_file_next[20][11] , \reg_file_next[20][10] ,
         \reg_file_next[20][9] , \reg_file_next[20][8] ,
         \reg_file_next[20][7] , \reg_file_next[20][6] ,
         \reg_file_next[20][5] , \reg_file_next[20][4] ,
         \reg_file_next[20][3] , \reg_file_next[20][2] ,
         \reg_file_next[20][1] , \reg_file_next[20][0] ,
         \reg_file_next[21][31] , \reg_file_next[21][30] ,
         \reg_file_next[21][29] , \reg_file_next[21][28] ,
         \reg_file_next[21][27] , \reg_file_next[21][26] ,
         \reg_file_next[21][25] , \reg_file_next[21][24] ,
         \reg_file_next[21][23] , \reg_file_next[21][22] ,
         \reg_file_next[21][21] , \reg_file_next[21][20] ,
         \reg_file_next[21][19] , \reg_file_next[21][18] ,
         \reg_file_next[21][17] , \reg_file_next[21][16] ,
         \reg_file_next[21][15] , \reg_file_next[21][14] ,
         \reg_file_next[21][13] , \reg_file_next[21][12] ,
         \reg_file_next[21][11] , \reg_file_next[21][10] ,
         \reg_file_next[21][9] , \reg_file_next[21][8] ,
         \reg_file_next[21][7] , \reg_file_next[21][6] ,
         \reg_file_next[21][5] , \reg_file_next[21][4] ,
         \reg_file_next[21][3] , \reg_file_next[21][2] ,
         \reg_file_next[21][1] , \reg_file_next[21][0] ,
         \reg_file_next[22][31] , \reg_file_next[22][30] ,
         \reg_file_next[22][29] , \reg_file_next[22][28] ,
         \reg_file_next[22][27] , \reg_file_next[22][26] ,
         \reg_file_next[22][25] , \reg_file_next[22][24] ,
         \reg_file_next[22][23] , \reg_file_next[22][22] ,
         \reg_file_next[22][21] , \reg_file_next[22][20] ,
         \reg_file_next[22][19] , \reg_file_next[22][18] ,
         \reg_file_next[22][17] , \reg_file_next[22][16] ,
         \reg_file_next[22][15] , \reg_file_next[22][14] ,
         \reg_file_next[22][13] , \reg_file_next[22][12] ,
         \reg_file_next[22][11] , \reg_file_next[22][10] ,
         \reg_file_next[22][9] , \reg_file_next[22][8] ,
         \reg_file_next[22][7] , \reg_file_next[22][6] ,
         \reg_file_next[22][5] , \reg_file_next[22][4] ,
         \reg_file_next[22][3] , \reg_file_next[22][2] ,
         \reg_file_next[22][1] , \reg_file_next[22][0] ,
         \reg_file_next[23][31] , \reg_file_next[23][30] ,
         \reg_file_next[23][29] , \reg_file_next[23][28] ,
         \reg_file_next[23][27] , \reg_file_next[23][26] ,
         \reg_file_next[23][25] , \reg_file_next[23][24] ,
         \reg_file_next[23][23] , \reg_file_next[23][22] ,
         \reg_file_next[23][21] , \reg_file_next[23][20] ,
         \reg_file_next[23][19] , \reg_file_next[23][18] ,
         \reg_file_next[23][17] , \reg_file_next[23][16] ,
         \reg_file_next[23][15] , \reg_file_next[23][14] ,
         \reg_file_next[23][13] , \reg_file_next[23][12] ,
         \reg_file_next[23][11] , \reg_file_next[23][10] ,
         \reg_file_next[23][9] , \reg_file_next[23][8] ,
         \reg_file_next[23][7] , \reg_file_next[23][6] ,
         \reg_file_next[23][5] , \reg_file_next[23][4] ,
         \reg_file_next[23][3] , \reg_file_next[23][2] ,
         \reg_file_next[23][1] , \reg_file_next[23][0] ,
         \reg_file_next[24][31] , \reg_file_next[24][30] ,
         \reg_file_next[24][29] , \reg_file_next[24][28] ,
         \reg_file_next[24][27] , \reg_file_next[24][26] ,
         \reg_file_next[24][25] , \reg_file_next[24][24] ,
         \reg_file_next[24][23] , \reg_file_next[24][22] ,
         \reg_file_next[24][21] , \reg_file_next[24][20] ,
         \reg_file_next[24][19] , \reg_file_next[24][18] ,
         \reg_file_next[24][17] , \reg_file_next[24][16] ,
         \reg_file_next[24][15] , \reg_file_next[24][14] ,
         \reg_file_next[24][13] , \reg_file_next[24][12] ,
         \reg_file_next[24][11] , \reg_file_next[24][10] ,
         \reg_file_next[24][9] , \reg_file_next[24][8] ,
         \reg_file_next[24][7] , \reg_file_next[24][6] ,
         \reg_file_next[24][5] , \reg_file_next[24][4] ,
         \reg_file_next[24][3] , \reg_file_next[24][2] ,
         \reg_file_next[24][1] , \reg_file_next[24][0] ,
         \reg_file_next[25][31] , \reg_file_next[25][30] ,
         \reg_file_next[25][29] , \reg_file_next[25][28] ,
         \reg_file_next[25][27] , \reg_file_next[25][26] ,
         \reg_file_next[25][25] , \reg_file_next[25][24] ,
         \reg_file_next[25][23] , \reg_file_next[25][22] ,
         \reg_file_next[25][21] , \reg_file_next[25][20] ,
         \reg_file_next[25][19] , \reg_file_next[25][18] ,
         \reg_file_next[25][17] , \reg_file_next[25][16] ,
         \reg_file_next[25][15] , \reg_file_next[25][14] ,
         \reg_file_next[25][13] , \reg_file_next[25][12] ,
         \reg_file_next[25][11] , \reg_file_next[25][10] ,
         \reg_file_next[25][9] , \reg_file_next[25][8] ,
         \reg_file_next[25][7] , \reg_file_next[25][6] ,
         \reg_file_next[25][5] , \reg_file_next[25][4] ,
         \reg_file_next[25][3] , \reg_file_next[25][2] ,
         \reg_file_next[25][1] , \reg_file_next[25][0] ,
         \reg_file_next[26][31] , \reg_file_next[26][30] ,
         \reg_file_next[26][29] , \reg_file_next[26][28] ,
         \reg_file_next[26][27] , \reg_file_next[26][26] ,
         \reg_file_next[26][25] , \reg_file_next[26][24] ,
         \reg_file_next[26][23] , \reg_file_next[26][22] ,
         \reg_file_next[26][21] , \reg_file_next[26][20] ,
         \reg_file_next[26][19] , \reg_file_next[26][18] ,
         \reg_file_next[26][17] , \reg_file_next[26][16] ,
         \reg_file_next[26][15] , \reg_file_next[26][14] ,
         \reg_file_next[26][13] , \reg_file_next[26][12] ,
         \reg_file_next[26][11] , \reg_file_next[26][10] ,
         \reg_file_next[26][9] , \reg_file_next[26][8] ,
         \reg_file_next[26][7] , \reg_file_next[26][6] ,
         \reg_file_next[26][5] , \reg_file_next[26][4] ,
         \reg_file_next[26][3] , \reg_file_next[26][2] ,
         \reg_file_next[26][1] , \reg_file_next[26][0] ,
         \reg_file_next[27][31] , \reg_file_next[27][30] ,
         \reg_file_next[27][29] , \reg_file_next[27][28] ,
         \reg_file_next[27][27] , \reg_file_next[27][26] ,
         \reg_file_next[27][25] , \reg_file_next[27][24] ,
         \reg_file_next[27][23] , \reg_file_next[27][22] ,
         \reg_file_next[27][21] , \reg_file_next[27][20] ,
         \reg_file_next[27][19] , \reg_file_next[27][18] ,
         \reg_file_next[27][17] , \reg_file_next[27][16] ,
         \reg_file_next[27][15] , \reg_file_next[27][14] ,
         \reg_file_next[27][13] , \reg_file_next[27][12] ,
         \reg_file_next[27][11] , \reg_file_next[27][10] ,
         \reg_file_next[27][9] , \reg_file_next[27][8] ,
         \reg_file_next[27][7] , \reg_file_next[27][6] ,
         \reg_file_next[27][5] , \reg_file_next[27][4] ,
         \reg_file_next[27][3] , \reg_file_next[27][2] ,
         \reg_file_next[27][1] , \reg_file_next[27][0] ,
         \reg_file_next[28][31] , \reg_file_next[28][30] ,
         \reg_file_next[28][29] , \reg_file_next[28][28] ,
         \reg_file_next[28][27] , \reg_file_next[28][26] ,
         \reg_file_next[28][25] , \reg_file_next[28][24] ,
         \reg_file_next[28][23] , \reg_file_next[28][22] ,
         \reg_file_next[28][21] , \reg_file_next[28][20] ,
         \reg_file_next[28][19] , \reg_file_next[28][18] ,
         \reg_file_next[28][17] , \reg_file_next[28][16] ,
         \reg_file_next[28][15] , \reg_file_next[28][14] ,
         \reg_file_next[28][13] , \reg_file_next[28][12] ,
         \reg_file_next[28][11] , \reg_file_next[28][10] ,
         \reg_file_next[28][9] , \reg_file_next[28][8] ,
         \reg_file_next[28][7] , \reg_file_next[28][6] ,
         \reg_file_next[28][5] , \reg_file_next[28][4] ,
         \reg_file_next[28][3] , \reg_file_next[28][2] ,
         \reg_file_next[28][1] , \reg_file_next[28][0] ,
         \reg_file_next[29][31] , \reg_file_next[29][30] ,
         \reg_file_next[29][29] , \reg_file_next[29][28] ,
         \reg_file_next[29][27] , \reg_file_next[29][26] ,
         \reg_file_next[29][25] , \reg_file_next[29][24] ,
         \reg_file_next[29][23] , \reg_file_next[29][22] ,
         \reg_file_next[29][21] , \reg_file_next[29][20] ,
         \reg_file_next[29][19] , \reg_file_next[29][18] ,
         \reg_file_next[29][17] , \reg_file_next[29][16] ,
         \reg_file_next[29][15] , \reg_file_next[29][14] ,
         \reg_file_next[29][13] , \reg_file_next[29][12] ,
         \reg_file_next[29][11] , \reg_file_next[29][10] ,
         \reg_file_next[29][9] , \reg_file_next[29][8] ,
         \reg_file_next[29][7] , \reg_file_next[29][6] ,
         \reg_file_next[29][5] , \reg_file_next[29][4] ,
         \reg_file_next[29][3] , \reg_file_next[29][2] ,
         \reg_file_next[29][1] , \reg_file_next[29][0] ,
         \reg_file_next[30][31] , \reg_file_next[30][30] ,
         \reg_file_next[30][29] , \reg_file_next[30][28] ,
         \reg_file_next[30][27] , \reg_file_next[30][26] ,
         \reg_file_next[30][25] , \reg_file_next[30][24] ,
         \reg_file_next[30][23] , \reg_file_next[30][22] ,
         \reg_file_next[30][21] , \reg_file_next[30][20] ,
         \reg_file_next[30][19] , \reg_file_next[30][18] ,
         \reg_file_next[30][17] , \reg_file_next[30][16] ,
         \reg_file_next[30][15] , \reg_file_next[30][14] ,
         \reg_file_next[30][13] , \reg_file_next[30][12] ,
         \reg_file_next[30][11] , \reg_file_next[30][10] ,
         \reg_file_next[30][9] , \reg_file_next[30][8] ,
         \reg_file_next[30][7] , \reg_file_next[30][6] ,
         \reg_file_next[30][5] , \reg_file_next[30][4] ,
         \reg_file_next[30][3] , \reg_file_next[30][2] ,
         \reg_file_next[30][1] , \reg_file_next[30][0] ,
         \reg_file_next[31][31] , \reg_file_next[31][30] ,
         \reg_file_next[31][29] , \reg_file_next[31][28] ,
         \reg_file_next[31][27] , \reg_file_next[31][26] ,
         \reg_file_next[31][25] , \reg_file_next[31][24] ,
         \reg_file_next[31][23] , \reg_file_next[31][22] ,
         \reg_file_next[31][21] , \reg_file_next[31][20] ,
         \reg_file_next[31][19] , \reg_file_next[31][18] ,
         \reg_file_next[31][17] , \reg_file_next[31][16] ,
         \reg_file_next[31][15] , \reg_file_next[31][14] ,
         \reg_file_next[31][13] , \reg_file_next[31][12] ,
         \reg_file_next[31][11] , \reg_file_next[31][10] ,
         \reg_file_next[31][9] , \reg_file_next[31][8] ,
         \reg_file_next[31][7] , \reg_file_next[31][6] ,
         \reg_file_next[31][5] , \reg_file_next[31][4] ,
         \reg_file_next[31][3] , \reg_file_next[31][2] ,
         \reg_file_next[31][1] , \reg_file_next[31][0] , Foward_C, Foward_D,
         N1140, \WB[0] , \EX[3] , n27, n28, n29, n30, n31, n70, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251;
  wire   [1:0] IR_addr;
  wire   [31:0] PC_plus4;
  wire   [31:0] PC_plus4Reg;
  wire   [31:0] InstReg;
  wire   [4:0] EX_Rt;
  wire   [2:0] EX_M;
  wire   [1:0] RegDST;
  wire   [1:0] Jump;
  wire   [2:0] ALUOp;
  wire   [2:0] WB_WB;
  wire   [4:0] WB_Rd;
  wire   [31:0] read_data1;
  wire   [31:0] read_data2;
  wire   [2:0] EX_WB;
  wire   [4:0] EX_Rd;
  wire   [31:0] after_C_MUX;
  wire   [31:0] aluresult;
  wire   [31:0] after_D_MUX;
  wire   [31:0] BranchAddr;
  wire   [2:0] M;
  wire   [2:0] WB_after_detect;
  wire   [2:0] MEM_after_detect;
  wire   [5:0] EX_after_detect;
  wire   [5:0] EX_reg;
  wire   [4:0] EX_Rs;
  wire   [31:0] EX_data1;
  wire   [31:0] EX_data2;
  wire   [31:0] EX_pcplus4;
  wire   [31:0] EX_signextend;
  wire   [3:0] ALUctrl;
  wire   [2:0] MEM_WB;
  wire   [4:0] MEM_Rd;
  wire   [1:0] Foward_A;
  wire   [1:0] Foward_B;
  wire   [31:0] after_A_mux;
  wire   [1:0] ALUOut_reg;
  wire   [31:0] after_B_mux;
  wire   [31:0] after_ALUSrc;
  wire   [31:0] MEM_pcplus4;
  wire   [31:0] WB_readdata;
  wire   [31:0] WB_ALUOut;
  wire   [31:0] WB_pcplus4;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign ICACHE_wdata[0] = 1'b0;
  assign ICACHE_wdata[1] = 1'b0;
  assign ICACHE_wdata[2] = 1'b0;
  assign ICACHE_wdata[3] = 1'b0;
  assign ICACHE_wdata[4] = 1'b0;
  assign ICACHE_wdata[5] = 1'b0;
  assign ICACHE_wdata[6] = 1'b0;
  assign ICACHE_wdata[7] = 1'b0;
  assign ICACHE_wdata[8] = 1'b0;
  assign ICACHE_wdata[9] = 1'b0;
  assign ICACHE_wdata[10] = 1'b0;
  assign ICACHE_wdata[11] = 1'b0;
  assign ICACHE_wdata[12] = 1'b0;
  assign ICACHE_wdata[13] = 1'b0;
  assign ICACHE_wdata[14] = 1'b0;
  assign ICACHE_wdata[15] = 1'b0;
  assign ICACHE_wdata[16] = 1'b0;
  assign ICACHE_wdata[17] = 1'b0;
  assign ICACHE_wdata[18] = 1'b0;
  assign ICACHE_wdata[19] = 1'b0;
  assign ICACHE_wdata[20] = 1'b0;
  assign ICACHE_wdata[21] = 1'b0;
  assign ICACHE_wdata[22] = 1'b0;
  assign ICACHE_wdata[23] = 1'b0;
  assign ICACHE_wdata[24] = 1'b0;
  assign ICACHE_wdata[25] = 1'b0;
  assign ICACHE_wdata[26] = 1'b0;
  assign ICACHE_wdata[27] = 1'b0;
  assign ICACHE_wdata[28] = 1'b0;
  assign ICACHE_wdata[29] = 1'b0;
  assign ICACHE_wdata[30] = 1'b0;
  assign ICACHE_wdata[31] = 1'b0;
  assign ICACHE_wen = 1'b0;
  assign ICACHE_ren = 1'b1;

  IFID IFID1 ( .IF_Flush(n2140), .clk(clk), .IFIDWrite(IFIDWrite), .PC_plus4(
        PC_plus4), .PC_plus4Reg(PC_plus4Reg), .Inst(ICACHE_rdata), .InstReg({
        InstReg[31:26], N72, N71, N70, N69, N68, N77, N76, N75, N74, N73, 
        InstReg[15:0]}), .stall_bothzero(n2209) );
  Hazard_detection hazard_detection ( .IDRegRS({N72, N71, N70, n2242, n2253}), 
        .IDRegRt({N77, N76, N75, n2210, n2224}), .EXRegRt(EX_Rt), .EXMemRead(
        EX_M[2]), .PCWrite(PCWrite), .IFIDWrite(IFIDWrite) );
  control control_unit ( .opcode(InstReg[31:26]), .rst_n(n2278), .Rs({N72, N71, 
        N70, n2242, n2253}), .Rt({N77, N76, N75, n2210, n2224}), .Rd(
        InstReg[15:11]), .RegDST(RegDST), .MemtoReg({SYNOPSYS_UNCONNECTED__0, 
        \MemtoReg[0] }), .Jump(Jump), .Branch(M[0]), .MemRead(M[2]), 
        .MemWrite(M[1]), .ALUSrc(\EX[3] ), .RegWrite(\WB[0] ), .ALUOp(ALUOp)
         );
  beq_foward beq_foward1 ( .RegWrite(EX_WB[0]), .instruction31_26(
        InstReg[31:26]), .instruction25_21({N72, N71, N70, n2242, n2253}), 
        .instruction20_16({N77, N76, N75, n2210, n2224}), .EX_Rd(EX_Rd), 
        .Foward_C(Foward_C), .Foward_D(Foward_D) );
  IDEX IDEX1 ( .clk(clk), .WB(WB_after_detect), .M(MEM_after_detect), .EX({
        WB_after_detect[2], EX_after_detect[4:0]}), .RegRs({N72, N71, N70, 
        n2242, n2253}), .RegRt({N77, N76, N75, n2210, n2224}), .RegRd(
        InstReg[15:11]), .data1(read_data1), .data2(read_data2), .sign_extend(
        {InstReg[15], InstReg[15], InstReg[15], InstReg[15], InstReg[15], 
        InstReg[15], InstReg[15], InstReg[15], InstReg[15], InstReg[15], 
        InstReg[15], InstReg[15], InstReg[15], InstReg[15], InstReg[15], 
        InstReg[15], InstReg[15:0]}), .PC_plus4Reg(PC_plus4Reg), .WB_reg(EX_WB), .M_reg(EX_M), .EX_reg(EX_reg), .RegRs_reg(EX_Rs), .RegRt_reg(EX_Rt), 
        .RegRd_reg(EX_Rd), .data1_reg(EX_data1), .data2_reg(EX_data2), 
        .EX_pcplus4(EX_pcplus4), .sign_extend_reg(EX_signextend), 
        .stall_bothzero(n2209) );
  ALUcontrol alucontrol ( .ALUctrl(ALUctrl), .ALUOp(EX_reg[2:0]), .func_field(
        EX_signextend[5:0]) );
  fowarding_unit fowarding_unit1 ( .ID_EX_Rs(EX_Rs), .ID_EX_Rt(EX_Rt), 
        .EX_MEM_RegWrite(MEM_WB[0]), .MEM_WB_RegWrite(WB_WB[0]), .EX_MEM_Rd(
        MEM_Rd), .MEM_WB_Rd(WB_Rd), .Foward_A(Foward_A), .Foward_B(Foward_B)
         );
  alu ALU ( .ALUin1(after_A_mux), .ALUin2(after_ALUSrc), .ALUctrl(ALUctrl), 
        .ALUresult(aluresult) );
  EXMEM EXMEM1 ( .clk(clk), .WB(EX_WB), .M(EX_M), .ALUOut(aluresult), .RegRD({
        n31, n30, n29, n28, n27}), .writedata(after_B_mux), .EX_pcplus4(
        EX_pcplus4), .WB_reg(MEM_WB), .M_reg({DCACHE_ren, DCACHE_wen, 
        SYNOPSYS_UNCONNECTED__1}), .ALUOut_reg({DCACHE_addr, ALUOut_reg}), 
        .RegRD_reg(MEM_Rd), .Writedata_reg(DCACHE_wdata), .stall_bothzero(
        n2209), .MEM_pcplus4(MEM_pcplus4) );
  MEMWB MEMWB1 ( .clk(clk), .WB(MEM_WB), .Memout(DCACHE_rdata), .ALUOut({
        DCACHE_addr, ALUOut_reg}), .RegRD(MEM_Rd), .MEM_pcplus4(MEM_pcplus4), 
        .WBreg(WB_WB), .Memreg(WB_readdata), .ALUreg(WB_ALUOut), .RegRDreg(
        WB_Rd), .stall_bothzero(n2209), .WB_pcplus4(WB_pcplus4) );
  MIPS_Pipeline_DW01_add_0 add_246 ( .A(PC_plus4Reg), .B({InstReg[15], 
        InstReg[15], InstReg[15], InstReg[15], InstReg[15], InstReg[15], 
        InstReg[15], InstReg[15], InstReg[15], InstReg[15], InstReg[15], 
        InstReg[15], InstReg[15], InstReg[15], InstReg[15:0], 1'b0, 1'b0}), 
        .CI(1'b0), .SUM(BranchAddr) );
  MIPS_Pipeline_DW01_cmp6_0 eq_233 ( .A(after_C_MUX), .B(after_D_MUX), .TC(
        1'b0), .EQ(N1140) );
  MIPS_Pipeline_DW01_add_1 add_156 ( .A({ICACHE_addr[29:1], n2130, IR_addr}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PC_plus4) );
  DFFRXL \IR_addr_reg[0]  ( .D(n1354), .CK(clk), .RN(n2285), .Q(IR_addr[0]), 
        .QN(n3251) );
  DFFRXL \IR_addr_reg[1]  ( .D(n1353), .CK(clk), .RN(n2285), .Q(IR_addr[1]), 
        .QN(n3250) );
  DFFRXL \reg_file_reg[0][31]  ( .D(n299), .CK(clk), .RN(n2282), .QN(n2129) );
  DFFRXL \reg_file_reg[0][30]  ( .D(n300), .CK(clk), .RN(n2271), .QN(n2128) );
  DFFRXL \reg_file_reg[0][29]  ( .D(n301), .CK(clk), .RN(n2271), .QN(n2127) );
  DFFRXL \reg_file_reg[0][28]  ( .D(n302), .CK(clk), .RN(n2272), .QN(n2126) );
  DFFRXL \reg_file_reg[0][27]  ( .D(n303), .CK(clk), .RN(n2272), .QN(n2125) );
  DFFRXL \reg_file_reg[0][26]  ( .D(n304), .CK(clk), .RN(n2273), .QN(n2124) );
  DFFRXL \reg_file_reg[0][25]  ( .D(n305), .CK(clk), .RN(n2273), .QN(n2123) );
  DFFRXL \reg_file_reg[0][24]  ( .D(n306), .CK(clk), .RN(n2283), .QN(n2122) );
  DFFRXL \reg_file_reg[0][23]  ( .D(n307), .CK(clk), .RN(n2284), .QN(n2121) );
  DFFRXL \reg_file_reg[0][22]  ( .D(n308), .CK(clk), .RN(n2274), .QN(n2120) );
  DFFRXL \reg_file_reg[0][21]  ( .D(n309), .CK(clk), .RN(n2274), .QN(n2119) );
  DFFRXL \reg_file_reg[0][20]  ( .D(n310), .CK(clk), .RN(n2279), .QN(n2118) );
  DFFRXL \reg_file_reg[0][19]  ( .D(n311), .CK(clk), .RN(n2275), .QN(n2117) );
  DFFRXL \reg_file_reg[0][18]  ( .D(n312), .CK(clk), .RN(n2284), .QN(n2116) );
  DFFRXL \reg_file_reg[0][17]  ( .D(n313), .CK(clk), .RN(n2275), .QN(n2115) );
  DFFRXL \reg_file_reg[0][16]  ( .D(n314), .CK(clk), .RN(n2276), .QN(n2114) );
  DFFRXL \reg_file_reg[0][15]  ( .D(n315), .CK(clk), .RN(n2276), .QN(n2113) );
  DFFRXL \reg_file_reg[0][14]  ( .D(n316), .CK(clk), .RN(n2277), .QN(n2112) );
  DFFRXL \reg_file_reg[0][13]  ( .D(n317), .CK(clk), .RN(n2277), .QN(n2111) );
  DFFRXL \reg_file_reg[0][12]  ( .D(n318), .CK(clk), .RN(n2278), .QN(n2110) );
  DFFRXL \reg_file_reg[0][11]  ( .D(n319), .CK(clk), .RN(n2278), .QN(n2109) );
  DFFRXL \reg_file_reg[0][10]  ( .D(n320), .CK(clk), .RN(n2279), .QN(n2108) );
  DFFRXL \reg_file_reg[0][9]  ( .D(n321), .CK(clk), .RN(n2279), .QN(n2107) );
  DFFRXL \reg_file_reg[0][8]  ( .D(n322), .CK(clk), .RN(n2280), .QN(n2106) );
  DFFRXL \reg_file_reg[0][7]  ( .D(n323), .CK(clk), .RN(n2281), .QN(n2105) );
  DFFRXL \reg_file_reg[0][6]  ( .D(n324), .CK(clk), .RN(n2281), .QN(n2104) );
  DFFRXL \reg_file_reg[0][5]  ( .D(n325), .CK(clk), .RN(n2284), .QN(n2103) );
  DFFRXL \reg_file_reg[0][4]  ( .D(n326), .CK(clk), .RN(n2284), .QN(n2102) );
  DFFRXL \reg_file_reg[0][3]  ( .D(n327), .CK(clk), .RN(n2284), .QN(n2101) );
  DFFRXL \reg_file_reg[0][2]  ( .D(n328), .CK(clk), .RN(n2282), .QN(n2100) );
  DFFRXL \reg_file_reg[0][1]  ( .D(n329), .CK(clk), .RN(n2284), .QN(n2099) );
  DFFRXL \reg_file_reg[0][0]  ( .D(n330), .CK(clk), .RN(n2284), .QN(n2098) );
  DFFRXL \reg_file_reg[1][31]  ( .D(n331), .CK(clk), .RN(n2279), .QN(n2097) );
  DFFRXL \reg_file_reg[1][30]  ( .D(n332), .CK(clk), .RN(n2271), .QN(n2096) );
  DFFRXL \reg_file_reg[1][29]  ( .D(n333), .CK(clk), .RN(n2271), .QN(n2095) );
  DFFRXL \reg_file_reg[1][28]  ( .D(n334), .CK(clk), .RN(n2272), .QN(n2094) );
  DFFRXL \reg_file_reg[1][27]  ( .D(n335), .CK(clk), .RN(n2272), .QN(n2093) );
  DFFRXL \reg_file_reg[1][26]  ( .D(n336), .CK(clk), .RN(n2273), .QN(n2092) );
  DFFRXL \reg_file_reg[1][25]  ( .D(n337), .CK(clk), .RN(n2273), .QN(n2091) );
  DFFRXL \reg_file_reg[1][24]  ( .D(n338), .CK(clk), .RN(n2282), .QN(n2090) );
  DFFRXL \reg_file_reg[1][23]  ( .D(n339), .CK(clk), .RN(n2278), .QN(n2089) );
  DFFRXL \reg_file_reg[1][22]  ( .D(n340), .CK(clk), .RN(n2274), .QN(n2088) );
  DFFRXL \reg_file_reg[1][21]  ( .D(n341), .CK(clk), .RN(n2274), .QN(n2087) );
  DFFRXL \reg_file_reg[1][20]  ( .D(n342), .CK(clk), .RN(n2271), .QN(n2086) );
  DFFRXL \reg_file_reg[1][19]  ( .D(n343), .CK(clk), .RN(n2275), .QN(n2085) );
  DFFRXL \reg_file_reg[1][18]  ( .D(n344), .CK(clk), .RN(n2284), .QN(n2084) );
  DFFRXL \reg_file_reg[1][17]  ( .D(n345), .CK(clk), .RN(n2275), .QN(n2083) );
  DFFRXL \reg_file_reg[1][16]  ( .D(n346), .CK(clk), .RN(n2276), .QN(n2082) );
  DFFRXL \reg_file_reg[1][15]  ( .D(n347), .CK(clk), .RN(n2276), .QN(n2081) );
  DFFRXL \reg_file_reg[1][14]  ( .D(n348), .CK(clk), .RN(n2277), .QN(n2080) );
  DFFRXL \reg_file_reg[1][13]  ( .D(n349), .CK(clk), .RN(n2277), .QN(n2079) );
  DFFRXL \reg_file_reg[1][12]  ( .D(n350), .CK(clk), .RN(n2278), .QN(n2078) );
  DFFRXL \reg_file_reg[1][11]  ( .D(n351), .CK(clk), .RN(n2278), .QN(n2077) );
  DFFRXL \reg_file_reg[1][10]  ( .D(n352), .CK(clk), .RN(n2279), .QN(n2076) );
  DFFRXL \reg_file_reg[1][9]  ( .D(n353), .CK(clk), .RN(n2279), .QN(n2075) );
  DFFRXL \reg_file_reg[1][8]  ( .D(n354), .CK(clk), .RN(n2280), .QN(n2074) );
  DFFRXL \reg_file_reg[1][7]  ( .D(n355), .CK(clk), .RN(n2281), .QN(n2073) );
  DFFRXL \reg_file_reg[1][6]  ( .D(n356), .CK(clk), .RN(n2281), .QN(n2072) );
  DFFRXL \reg_file_reg[1][5]  ( .D(n357), .CK(clk), .RN(n2284), .QN(n2071) );
  DFFRXL \reg_file_reg[1][4]  ( .D(n358), .CK(clk), .RN(n2284), .QN(n2070) );
  DFFRXL \reg_file_reg[1][3]  ( .D(n359), .CK(clk), .RN(n2284), .QN(n2069) );
  DFFRXL \reg_file_reg[1][2]  ( .D(n360), .CK(clk), .RN(n2282), .QN(n2068) );
  DFFRXL \reg_file_reg[1][1]  ( .D(n361), .CK(clk), .RN(n2284), .QN(n2067) );
  DFFRXL \reg_file_reg[1][0]  ( .D(n362), .CK(clk), .RN(n2284), .QN(n2066) );
  DFFRXL \reg_file_reg[2][31]  ( .D(n363), .CK(clk), .RN(n2274), .QN(n2065) );
  DFFRXL \reg_file_reg[2][30]  ( .D(n364), .CK(clk), .RN(n2277), .QN(n2064) );
  DFFRXL \reg_file_reg[2][29]  ( .D(n365), .CK(clk), .RN(n2271), .QN(n2063) );
  DFFRXL \reg_file_reg[2][28]  ( .D(n366), .CK(clk), .RN(n2272), .QN(n2062) );
  DFFRXL \reg_file_reg[2][27]  ( .D(n367), .CK(clk), .RN(n2272), .QN(n2061) );
  DFFRXL \reg_file_reg[2][26]  ( .D(n368), .CK(clk), .RN(n2273), .QN(n2060) );
  DFFRXL \reg_file_reg[2][25]  ( .D(n369), .CK(clk), .RN(n2273), .QN(n2059) );
  DFFRXL \reg_file_reg[2][24]  ( .D(n370), .CK(clk), .RN(n2279), .QN(n2058) );
  DFFRXL \reg_file_reg[2][23]  ( .D(n371), .CK(clk), .RN(n2271), .QN(n2057) );
  DFFRXL \reg_file_reg[2][22]  ( .D(n372), .CK(clk), .RN(n2274), .QN(n2056) );
  DFFRXL \reg_file_reg[2][21]  ( .D(n373), .CK(clk), .RN(n2274), .QN(n2055) );
  DFFRXL \reg_file_reg[2][20]  ( .D(n374), .CK(clk), .RN(n2274), .QN(n2054) );
  DFFRXL \reg_file_reg[2][19]  ( .D(n375), .CK(clk), .RN(n2275), .QN(n2053) );
  DFFRXL \reg_file_reg[2][18]  ( .D(n376), .CK(clk), .RN(n2284), .QN(n2052) );
  DFFRXL \reg_file_reg[2][17]  ( .D(n377), .CK(clk), .RN(n2275), .QN(n2051) );
  DFFRXL \reg_file_reg[2][16]  ( .D(n378), .CK(clk), .RN(n2276), .QN(n2050) );
  DFFRXL \reg_file_reg[2][15]  ( .D(n379), .CK(clk), .RN(n2276), .QN(n2049) );
  DFFRXL \reg_file_reg[2][14]  ( .D(n380), .CK(clk), .RN(n2277), .QN(n2048) );
  DFFRXL \reg_file_reg[2][13]  ( .D(n381), .CK(clk), .RN(n2277), .QN(n2047) );
  DFFRXL \reg_file_reg[2][12]  ( .D(n382), .CK(clk), .RN(n2278), .QN(n2046) );
  DFFRXL \reg_file_reg[2][11]  ( .D(n383), .CK(clk), .RN(n2278), .QN(n2045) );
  DFFRXL \reg_file_reg[2][10]  ( .D(n384), .CK(clk), .RN(n2279), .QN(n2044) );
  DFFRXL \reg_file_reg[2][9]  ( .D(n385), .CK(clk), .RN(n2279), .QN(n2043) );
  DFFRXL \reg_file_reg[2][8]  ( .D(n386), .CK(clk), .RN(n2280), .QN(n2042) );
  DFFRXL \reg_file_reg[2][7]  ( .D(n387), .CK(clk), .RN(n2281), .QN(n2041) );
  DFFRXL \reg_file_reg[2][6]  ( .D(n388), .CK(clk), .RN(n2281), .QN(n2040) );
  DFFRXL \reg_file_reg[2][5]  ( .D(n389), .CK(clk), .RN(n2284), .QN(n2039) );
  DFFRXL \reg_file_reg[2][4]  ( .D(n390), .CK(clk), .RN(n2284), .QN(n2038) );
  DFFRXL \reg_file_reg[2][3]  ( .D(n391), .CK(clk), .RN(n2284), .QN(n2037) );
  DFFRXL \reg_file_reg[2][2]  ( .D(n392), .CK(clk), .RN(n2282), .QN(n2036) );
  DFFRXL \reg_file_reg[2][1]  ( .D(n393), .CK(clk), .RN(n2284), .QN(n2035) );
  DFFRXL \reg_file_reg[2][0]  ( .D(n394), .CK(clk), .RN(n2284), .QN(n2034) );
  DFFRXL \reg_file_reg[3][31]  ( .D(n395), .CK(clk), .RN(n2273), .QN(n2033) );
  DFFRXL \reg_file_reg[3][30]  ( .D(n396), .CK(clk), .RN(n2272), .QN(n2032) );
  DFFRXL \reg_file_reg[3][29]  ( .D(n397), .CK(clk), .RN(n2271), .QN(n2031) );
  DFFRXL \reg_file_reg[3][28]  ( .D(n398), .CK(clk), .RN(n2272), .QN(n2030) );
  DFFRXL \reg_file_reg[3][27]  ( .D(n399), .CK(clk), .RN(n2272), .QN(n2029) );
  DFFRXL \reg_file_reg[3][26]  ( .D(n400), .CK(clk), .RN(n2273), .QN(n2028) );
  DFFRXL \reg_file_reg[3][25]  ( .D(n401), .CK(clk), .RN(n2273), .QN(n2027) );
  DFFRXL \reg_file_reg[3][24]  ( .D(n402), .CK(clk), .RN(n2274), .QN(n2026) );
  DFFRXL \reg_file_reg[3][23]  ( .D(n403), .CK(clk), .RN(n2277), .QN(n2025) );
  DFFRXL \reg_file_reg[3][22]  ( .D(n404), .CK(clk), .RN(n2274), .QN(n2024) );
  DFFRXL \reg_file_reg[3][21]  ( .D(n405), .CK(clk), .RN(n2274), .QN(n2023) );
  DFFRXL \reg_file_reg[3][20]  ( .D(n406), .CK(clk), .RN(n2277), .QN(n2022) );
  DFFRXL \reg_file_reg[3][19]  ( .D(n407), .CK(clk), .RN(n2275), .QN(n2021) );
  DFFRXL \reg_file_reg[3][18]  ( .D(n408), .CK(clk), .RN(n2284), .QN(n2020) );
  DFFRXL \reg_file_reg[3][17]  ( .D(n409), .CK(clk), .RN(n2275), .QN(n2019) );
  DFFRXL \reg_file_reg[3][16]  ( .D(n410), .CK(clk), .RN(n2276), .QN(n2018) );
  DFFRXL \reg_file_reg[3][15]  ( .D(n411), .CK(clk), .RN(n2276), .QN(n2017) );
  DFFRXL \reg_file_reg[3][14]  ( .D(n412), .CK(clk), .RN(n2277), .QN(n2016) );
  DFFRXL \reg_file_reg[3][13]  ( .D(n413), .CK(clk), .RN(n2277), .QN(n2015) );
  DFFRXL \reg_file_reg[3][12]  ( .D(n414), .CK(clk), .RN(n2278), .QN(n2014) );
  DFFRXL \reg_file_reg[3][11]  ( .D(n415), .CK(clk), .RN(n2278), .QN(n2013) );
  DFFRXL \reg_file_reg[3][10]  ( .D(n416), .CK(clk), .RN(n2279), .QN(n2012) );
  DFFRXL \reg_file_reg[3][9]  ( .D(n417), .CK(clk), .RN(n2279), .QN(n2011) );
  DFFRXL \reg_file_reg[3][8]  ( .D(n418), .CK(clk), .RN(n2280), .QN(n2010) );
  DFFRXL \reg_file_reg[3][7]  ( .D(n419), .CK(clk), .RN(n2281), .QN(n2009) );
  DFFRXL \reg_file_reg[3][6]  ( .D(n420), .CK(clk), .RN(n2281), .QN(n2008) );
  DFFRXL \reg_file_reg[3][5]  ( .D(n421), .CK(clk), .RN(n2284), .QN(n2007) );
  DFFRXL \reg_file_reg[3][4]  ( .D(n422), .CK(clk), .RN(n2284), .QN(n2006) );
  DFFRXL \reg_file_reg[3][3]  ( .D(n423), .CK(clk), .RN(n2284), .QN(n2005) );
  DFFRXL \reg_file_reg[3][2]  ( .D(n424), .CK(clk), .RN(n2282), .QN(n2004) );
  DFFRXL \reg_file_reg[3][1]  ( .D(n425), .CK(clk), .RN(n2284), .QN(n2003) );
  DFFRXL \reg_file_reg[3][0]  ( .D(n426), .CK(clk), .RN(n2284), .QN(n2002) );
  DFFRXL \reg_file_reg[4][31]  ( .D(n427), .CK(clk), .RN(n2276), .QN(n2001) );
  DFFRXL \reg_file_reg[4][30]  ( .D(n428), .CK(clk), .RN(n2274), .QN(n2000) );
  DFFRXL \reg_file_reg[4][29]  ( .D(n429), .CK(clk), .RN(n2271), .QN(n1999) );
  DFFRXL \reg_file_reg[4][28]  ( .D(n430), .CK(clk), .RN(n2272), .QN(n1998) );
  DFFRXL \reg_file_reg[4][27]  ( .D(n431), .CK(clk), .RN(n2272), .QN(n1997) );
  DFFRXL \reg_file_reg[4][26]  ( .D(n432), .CK(clk), .RN(n2273), .QN(n1996) );
  DFFRXL \reg_file_reg[4][25]  ( .D(n433), .CK(clk), .RN(n2273), .QN(n1995) );
  DFFRXL \reg_file_reg[4][24]  ( .D(n434), .CK(clk), .RN(n2273), .QN(n1994) );
  DFFRXL \reg_file_reg[4][23]  ( .D(n435), .CK(clk), .RN(n2272), .QN(n1993) );
  DFFRXL \reg_file_reg[4][22]  ( .D(n436), .CK(clk), .RN(n2274), .QN(n1992) );
  DFFRXL \reg_file_reg[4][21]  ( .D(n437), .CK(clk), .RN(n2274), .QN(n1991) );
  DFFRXL \reg_file_reg[4][20]  ( .D(n438), .CK(clk), .RN(n2273), .QN(n1990) );
  DFFRXL \reg_file_reg[4][19]  ( .D(n439), .CK(clk), .RN(n2272), .QN(n1989) );
  DFFRXL \reg_file_reg[4][18]  ( .D(n440), .CK(clk), .RN(n2284), .QN(n1988) );
  DFFRXL \reg_file_reg[4][17]  ( .D(n441), .CK(clk), .RN(n2275), .QN(n1987) );
  DFFRXL \reg_file_reg[4][16]  ( .D(n442), .CK(clk), .RN(n2276), .QN(n1986) );
  DFFRXL \reg_file_reg[4][15]  ( .D(n443), .CK(clk), .RN(n2276), .QN(n1985) );
  DFFRXL \reg_file_reg[4][14]  ( .D(n444), .CK(clk), .RN(n2277), .QN(n1984) );
  DFFRXL \reg_file_reg[4][13]  ( .D(n445), .CK(clk), .RN(n2277), .QN(n1983) );
  DFFRXL \reg_file_reg[4][12]  ( .D(n446), .CK(clk), .RN(n2278), .QN(n1982) );
  DFFRXL \reg_file_reg[4][11]  ( .D(n447), .CK(clk), .RN(n2278), .QN(n1981) );
  DFFRXL \reg_file_reg[4][10]  ( .D(n448), .CK(clk), .RN(n2279), .QN(n1980) );
  DFFRXL \reg_file_reg[4][9]  ( .D(n449), .CK(clk), .RN(n2279), .QN(n1979) );
  DFFRXL \reg_file_reg[4][8]  ( .D(n450), .CK(clk), .RN(n2280), .QN(n1978) );
  DFFRXL \reg_file_reg[4][7]  ( .D(n451), .CK(clk), .RN(n2281), .QN(n1977) );
  DFFRXL \reg_file_reg[4][6]  ( .D(n452), .CK(clk), .RN(n2281), .QN(n1976) );
  DFFRXL \reg_file_reg[4][5]  ( .D(n453), .CK(clk), .RN(n2284), .QN(n1975) );
  DFFRXL \reg_file_reg[4][4]  ( .D(n454), .CK(clk), .RN(n2284), .QN(n1974) );
  DFFRXL \reg_file_reg[4][3]  ( .D(n455), .CK(clk), .RN(n2284), .QN(n1973) );
  DFFRXL \reg_file_reg[4][2]  ( .D(n456), .CK(clk), .RN(n2282), .QN(n1972) );
  DFFRXL \reg_file_reg[4][1]  ( .D(n457), .CK(clk), .RN(n2284), .QN(n1971) );
  DFFRXL \reg_file_reg[4][0]  ( .D(n458), .CK(clk), .RN(n2284), .QN(n1970) );
  DFFRXL \reg_file_reg[5][31]  ( .D(n459), .CK(clk), .RN(n2275), .QN(n1969) );
  DFFRXL \reg_file_reg[5][30]  ( .D(n460), .CK(clk), .RN(n2280), .QN(n1968) );
  DFFRXL \reg_file_reg[5][29]  ( .D(n461), .CK(clk), .RN(n2271), .QN(n1967) );
  DFFRXL \reg_file_reg[5][28]  ( .D(n462), .CK(clk), .RN(n2272), .QN(n1966) );
  DFFRXL \reg_file_reg[5][27]  ( .D(n463), .CK(clk), .RN(n2272), .QN(n1965) );
  DFFRXL \reg_file_reg[5][26]  ( .D(n464), .CK(clk), .RN(n2273), .QN(n1964) );
  DFFRXL \reg_file_reg[5][25]  ( .D(n465), .CK(clk), .RN(n2273), .QN(n1963) );
  DFFRXL \reg_file_reg[5][24]  ( .D(n466), .CK(clk), .RN(n2276), .QN(n1962) );
  DFFRXL \reg_file_reg[5][23]  ( .D(n467), .CK(clk), .RN(n2272), .QN(n1961) );
  DFFRXL \reg_file_reg[5][22]  ( .D(n468), .CK(clk), .RN(n2274), .QN(n1960) );
  DFFRXL \reg_file_reg[5][21]  ( .D(n469), .CK(clk), .RN(n2274), .QN(n1959) );
  DFFRXL \reg_file_reg[5][20]  ( .D(n470), .CK(clk), .RN(n2281), .QN(n1958) );
  DFFRXL \reg_file_reg[5][19]  ( .D(n471), .CK(clk), .RN(n2276), .QN(n1957) );
  DFFRXL \reg_file_reg[5][18]  ( .D(n472), .CK(clk), .RN(n2284), .QN(n1956) );
  DFFRXL \reg_file_reg[5][17]  ( .D(n473), .CK(clk), .RN(n2275), .QN(n1955) );
  DFFRXL \reg_file_reg[5][16]  ( .D(n474), .CK(clk), .RN(n2276), .QN(n1954) );
  DFFRXL \reg_file_reg[5][15]  ( .D(n475), .CK(clk), .RN(n2276), .QN(n1953) );
  DFFRXL \reg_file_reg[5][14]  ( .D(n476), .CK(clk), .RN(n2277), .QN(n1952) );
  DFFRXL \reg_file_reg[5][13]  ( .D(n477), .CK(clk), .RN(n2277), .QN(n1951) );
  DFFRXL \reg_file_reg[5][12]  ( .D(n478), .CK(clk), .RN(n2278), .QN(n1950) );
  DFFRXL \reg_file_reg[5][11]  ( .D(n479), .CK(clk), .RN(n2278), .QN(n1949) );
  DFFRXL \reg_file_reg[5][10]  ( .D(n480), .CK(clk), .RN(n2279), .QN(n1948) );
  DFFRXL \reg_file_reg[5][9]  ( .D(n481), .CK(clk), .RN(n2279), .QN(n1947) );
  DFFRXL \reg_file_reg[5][8]  ( .D(n482), .CK(clk), .RN(n2280), .QN(n1946) );
  DFFRXL \reg_file_reg[5][7]  ( .D(n483), .CK(clk), .RN(n2281), .QN(n1945) );
  DFFRXL \reg_file_reg[5][6]  ( .D(n484), .CK(clk), .RN(n2281), .QN(n1944) );
  DFFRXL \reg_file_reg[5][5]  ( .D(n485), .CK(clk), .RN(n2284), .QN(n1943) );
  DFFRXL \reg_file_reg[5][4]  ( .D(n486), .CK(clk), .RN(n2284), .QN(n1942) );
  DFFRXL \reg_file_reg[5][3]  ( .D(n487), .CK(clk), .RN(n2284), .QN(n1941) );
  DFFRXL \reg_file_reg[5][2]  ( .D(n488), .CK(clk), .RN(n2282), .QN(n1940) );
  DFFRXL \reg_file_reg[5][1]  ( .D(n489), .CK(clk), .RN(n2284), .QN(n1939) );
  DFFRXL \reg_file_reg[5][0]  ( .D(n490), .CK(clk), .RN(n2284), .QN(n1938) );
  DFFRXL \reg_file_reg[6][31]  ( .D(n491), .CK(clk), .RN(n2281), .QN(n1937) );
  DFFRXL \reg_file_reg[6][30]  ( .D(n492), .CK(clk), .RN(n2281), .QN(n1936) );
  DFFRXL \reg_file_reg[6][29]  ( .D(n493), .CK(clk), .RN(n2271), .QN(n1935) );
  DFFRXL \reg_file_reg[6][28]  ( .D(n494), .CK(clk), .RN(n2272), .QN(n1934) );
  DFFRXL \reg_file_reg[6][27]  ( .D(n495), .CK(clk), .RN(n2272), .QN(n1933) );
  DFFRXL \reg_file_reg[6][26]  ( .D(n496), .CK(clk), .RN(n2273), .QN(n1932) );
  DFFRXL \reg_file_reg[6][25]  ( .D(n497), .CK(clk), .RN(n2273), .QN(n1931) );
  DFFRXL \reg_file_reg[6][24]  ( .D(n498), .CK(clk), .RN(n2275), .QN(n1930) );
  DFFRXL \reg_file_reg[6][23]  ( .D(n499), .CK(clk), .RN(n2280), .QN(n1929) );
  DFFRXL \reg_file_reg[6][22]  ( .D(n500), .CK(clk), .RN(n2274), .QN(n1928) );
  DFFRXL \reg_file_reg[6][21]  ( .D(n501), .CK(clk), .RN(n2274), .QN(n1927) );
  DFFRXL \reg_file_reg[6][20]  ( .D(n502), .CK(clk), .RN(n2275), .QN(n1926) );
  DFFRXL \reg_file_reg[6][19]  ( .D(n503), .CK(clk), .RN(n2280), .QN(n1925) );
  DFFRXL \reg_file_reg[6][18]  ( .D(n504), .CK(clk), .RN(n2284), .QN(n1924) );
  DFFRXL \reg_file_reg[6][17]  ( .D(n505), .CK(clk), .RN(n2275), .QN(n1923) );
  DFFRXL \reg_file_reg[6][16]  ( .D(n506), .CK(clk), .RN(n2276), .QN(n1922) );
  DFFRXL \reg_file_reg[6][15]  ( .D(n507), .CK(clk), .RN(n2276), .QN(n1921) );
  DFFRXL \reg_file_reg[6][14]  ( .D(n508), .CK(clk), .RN(n2277), .QN(n1920) );
  DFFRXL \reg_file_reg[6][13]  ( .D(n509), .CK(clk), .RN(n2277), .QN(n1919) );
  DFFRXL \reg_file_reg[6][12]  ( .D(n510), .CK(clk), .RN(n2278), .QN(n1918) );
  DFFRXL \reg_file_reg[6][11]  ( .D(n511), .CK(clk), .RN(n2278), .QN(n1917) );
  DFFRXL \reg_file_reg[6][10]  ( .D(n512), .CK(clk), .RN(n2279), .QN(n1916) );
  DFFRXL \reg_file_reg[6][9]  ( .D(n513), .CK(clk), .RN(n2279), .QN(n1915) );
  DFFRXL \reg_file_reg[6][8]  ( .D(n514), .CK(clk), .RN(n2280), .QN(n1914) );
  DFFRXL \reg_file_reg[6][7]  ( .D(n515), .CK(clk), .RN(n2280), .QN(n1913) );
  DFFRXL \reg_file_reg[6][6]  ( .D(n516), .CK(clk), .RN(n2281), .QN(n1912) );
  DFFRXL \reg_file_reg[6][5]  ( .D(n517), .CK(clk), .RN(n2284), .QN(n1911) );
  DFFRXL \reg_file_reg[6][4]  ( .D(n518), .CK(clk), .RN(n2284), .QN(n1910) );
  DFFRXL \reg_file_reg[6][3]  ( .D(n519), .CK(clk), .RN(n2284), .QN(n1909) );
  DFFRXL \reg_file_reg[6][2]  ( .D(n520), .CK(clk), .RN(n2282), .QN(n1908) );
  DFFRXL \reg_file_reg[6][1]  ( .D(n521), .CK(clk), .RN(n2284), .QN(n1907) );
  DFFRXL \reg_file_reg[6][0]  ( .D(n522), .CK(clk), .RN(n2284), .QN(n1906) );
  DFFRXL \reg_file_reg[7][31]  ( .D(n523), .CK(clk), .RN(n2283), .QN(n1905) );
  DFFRXL \reg_file_reg[7][30]  ( .D(n524), .CK(clk), .RN(n2284), .QN(n1904) );
  DFFRXL \reg_file_reg[7][29]  ( .D(n525), .CK(clk), .RN(n2271), .QN(n1903) );
  DFFRXL \reg_file_reg[7][28]  ( .D(n526), .CK(clk), .RN(n2271), .QN(n1902) );
  DFFRXL \reg_file_reg[7][27]  ( .D(n527), .CK(clk), .RN(n2272), .QN(n1901) );
  DFFRXL \reg_file_reg[7][26]  ( .D(n528), .CK(clk), .RN(n2273), .QN(n1900) );
  DFFRXL \reg_file_reg[7][25]  ( .D(n529), .CK(clk), .RN(n2273), .QN(n1899) );
  DFFRXL \reg_file_reg[7][24]  ( .D(n530), .CK(clk), .RN(n2281), .QN(n1898) );
  DFFRXL \reg_file_reg[7][23]  ( .D(n531), .CK(clk), .RN(n2283), .QN(n1897) );
  DFFRXL \reg_file_reg[7][22]  ( .D(n532), .CK(clk), .RN(n2274), .QN(n1896) );
  DFFRXL \reg_file_reg[7][21]  ( .D(n533), .CK(clk), .RN(n2274), .QN(n1895) );
  DFFRXL \reg_file_reg[7][20]  ( .D(n534), .CK(clk), .RN(n2283), .QN(n1894) );
  DFFRXL \reg_file_reg[7][19]  ( .D(n535), .CK(clk), .RN(n2284), .QN(n1893) );
  DFFRXL \reg_file_reg[7][18]  ( .D(n536), .CK(clk), .RN(n2284), .QN(n1892) );
  DFFRXL \reg_file_reg[7][17]  ( .D(n537), .CK(clk), .RN(n2275), .QN(n1891) );
  DFFRXL \reg_file_reg[7][16]  ( .D(n538), .CK(clk), .RN(n2276), .QN(n1890) );
  DFFRXL \reg_file_reg[7][15]  ( .D(n539), .CK(clk), .RN(n2276), .QN(n1889) );
  DFFRXL \reg_file_reg[7][14]  ( .D(n540), .CK(clk), .RN(n2277), .QN(n1888) );
  DFFRXL \reg_file_reg[7][13]  ( .D(n541), .CK(clk), .RN(n2277), .QN(n1887) );
  DFFRXL \reg_file_reg[7][12]  ( .D(n542), .CK(clk), .RN(n2278), .QN(n1886) );
  DFFRXL \reg_file_reg[7][11]  ( .D(n543), .CK(clk), .RN(n2278), .QN(n1885) );
  DFFRXL \reg_file_reg[7][10]  ( .D(n544), .CK(clk), .RN(n2279), .QN(n1884) );
  DFFRXL \reg_file_reg[7][9]  ( .D(n545), .CK(clk), .RN(n2279), .QN(n1883) );
  DFFRXL \reg_file_reg[7][8]  ( .D(n546), .CK(clk), .RN(n2280), .QN(n1882) );
  DFFRXL \reg_file_reg[7][7]  ( .D(n547), .CK(clk), .RN(n2280), .QN(n1881) );
  DFFRXL \reg_file_reg[7][6]  ( .D(n548), .CK(clk), .RN(n2281), .QN(n1880) );
  DFFRXL \reg_file_reg[7][5]  ( .D(n549), .CK(clk), .RN(n2284), .QN(n1879) );
  DFFRXL \reg_file_reg[7][4]  ( .D(n550), .CK(clk), .RN(n2284), .QN(n1878) );
  DFFRXL \reg_file_reg[7][3]  ( .D(n551), .CK(clk), .RN(n2283), .QN(n1877) );
  DFFRXL \reg_file_reg[7][2]  ( .D(n552), .CK(clk), .RN(n2282), .QN(n1876) );
  DFFRXL \reg_file_reg[7][1]  ( .D(n553), .CK(clk), .RN(n2283), .QN(n1875) );
  DFFRXL \reg_file_reg[7][0]  ( .D(n554), .CK(clk), .RN(n2283), .QN(n1874) );
  DFFRXL \reg_file_reg[8][31]  ( .D(n555), .CK(clk), .RN(n2278), .QN(n1873) );
  DFFRXL \reg_file_reg[8][30]  ( .D(n556), .CK(clk), .RN(n2282), .QN(n1872) );
  DFFRXL \reg_file_reg[8][29]  ( .D(n557), .CK(clk), .RN(n2271), .QN(n1871) );
  DFFRXL \reg_file_reg[8][28]  ( .D(n558), .CK(clk), .RN(n2271), .QN(n1870) );
  DFFRXL \reg_file_reg[8][27]  ( .D(n559), .CK(clk), .RN(n2272), .QN(n1869) );
  DFFRXL \reg_file_reg[8][26]  ( .D(n560), .CK(clk), .RN(n2273), .QN(n1868) );
  DFFRXL \reg_file_reg[8][25]  ( .D(n561), .CK(clk), .RN(n2273), .QN(n1867) );
  DFFRXL \reg_file_reg[8][24]  ( .D(n562), .CK(clk), .RN(n2284), .QN(n1866) );
  DFFRXL \reg_file_reg[8][23]  ( .D(n563), .CK(clk), .RN(n2282), .QN(n1865) );
  DFFRXL \reg_file_reg[8][22]  ( .D(n564), .CK(clk), .RN(n2274), .QN(n1864) );
  DFFRXL \reg_file_reg[8][21]  ( .D(n565), .CK(clk), .RN(n2274), .QN(n1863) );
  DFFRXL \reg_file_reg[8][20]  ( .D(n566), .CK(clk), .RN(n2282), .QN(n1862) );
  DFFRXL \reg_file_reg[8][19]  ( .D(n567), .CK(clk), .RN(n2278), .QN(n1861) );
  DFFRXL \reg_file_reg[8][18]  ( .D(n568), .CK(clk), .RN(n2285), .QN(n1860) );
  DFFRXL \reg_file_reg[8][17]  ( .D(n569), .CK(clk), .RN(n2275), .QN(n1859) );
  DFFRXL \reg_file_reg[8][16]  ( .D(n570), .CK(clk), .RN(n2276), .QN(n1858) );
  DFFRXL \reg_file_reg[8][15]  ( .D(n571), .CK(clk), .RN(n2276), .QN(n1857) );
  DFFRXL \reg_file_reg[8][14]  ( .D(n572), .CK(clk), .RN(n2277), .QN(n1856) );
  DFFRXL \reg_file_reg[8][13]  ( .D(n573), .CK(clk), .RN(n2277), .QN(n1855) );
  DFFRXL \reg_file_reg[8][12]  ( .D(n574), .CK(clk), .RN(n2278), .QN(n1854) );
  DFFRXL \reg_file_reg[8][11]  ( .D(n575), .CK(clk), .RN(n2278), .QN(n1853) );
  DFFRXL \reg_file_reg[8][10]  ( .D(n576), .CK(clk), .RN(n2279), .QN(n1852) );
  DFFRXL \reg_file_reg[8][9]  ( .D(n577), .CK(clk), .RN(n2279), .QN(n1851) );
  DFFRXL \reg_file_reg[8][8]  ( .D(n578), .CK(clk), .RN(n2280), .QN(n1850) );
  DFFRXL \reg_file_reg[8][7]  ( .D(n579), .CK(clk), .RN(n2280), .QN(n1849) );
  DFFRXL \reg_file_reg[8][6]  ( .D(n580), .CK(clk), .RN(n2281), .QN(n1848) );
  DFFRXL \reg_file_reg[8][5]  ( .D(n581), .CK(clk), .RN(n2285), .QN(n1847) );
  DFFRXL \reg_file_reg[8][4]  ( .D(n582), .CK(clk), .RN(n2285), .QN(n1846) );
  DFFRXL \reg_file_reg[8][3]  ( .D(n583), .CK(clk), .RN(n2285), .QN(n1845) );
  DFFRXL \reg_file_reg[8][2]  ( .D(n584), .CK(clk), .RN(n2282), .QN(n1844) );
  DFFRXL \reg_file_reg[8][1]  ( .D(n585), .CK(clk), .RN(n2285), .QN(n1843) );
  DFFRXL \reg_file_reg[8][0]  ( .D(n586), .CK(clk), .RN(n2285), .QN(n1842) );
  DFFRXL \reg_file_reg[9][31]  ( .D(n587), .CK(clk), .RN(n2279), .QN(n1841) );
  DFFRXL \reg_file_reg[9][30]  ( .D(n588), .CK(clk), .RN(n2271), .QN(n1840) );
  DFFRXL \reg_file_reg[9][29]  ( .D(n589), .CK(clk), .RN(n2271), .QN(n1839) );
  DFFRXL \reg_file_reg[9][28]  ( .D(n590), .CK(clk), .RN(n2271), .QN(n1838) );
  DFFRXL \reg_file_reg[9][27]  ( .D(n591), .CK(clk), .RN(n2272), .QN(n1837) );
  DFFRXL \reg_file_reg[9][26]  ( .D(n592), .CK(clk), .RN(n2273), .QN(n1836) );
  DFFRXL \reg_file_reg[9][25]  ( .D(n593), .CK(clk), .RN(n2273), .QN(n1835) );
  DFFRXL \reg_file_reg[9][24]  ( .D(n594), .CK(clk), .RN(n2278), .QN(n1834) );
  DFFRXL \reg_file_reg[9][23]  ( .D(n595), .CK(clk), .RN(n2279), .QN(n1833) );
  DFFRXL \reg_file_reg[9][22]  ( .D(n596), .CK(clk), .RN(n2274), .QN(n1832) );
  DFFRXL \reg_file_reg[9][21]  ( .D(n597), .CK(clk), .RN(n2274), .QN(n1831) );
  DFFRXL \reg_file_reg[9][20]  ( .D(n598), .CK(clk), .RN(n2279), .QN(n1830) );
  DFFRXL \reg_file_reg[9][19]  ( .D(n599), .CK(clk), .RN(n2271), .QN(n1829) );
  DFFRXL \reg_file_reg[9][18]  ( .D(n600), .CK(clk), .RN(n2285), .QN(n1828) );
  DFFRXL \reg_file_reg[9][17]  ( .D(n601), .CK(clk), .RN(n2275), .QN(n1827) );
  DFFRXL \reg_file_reg[9][16]  ( .D(n602), .CK(clk), .RN(n2276), .QN(n1826) );
  DFFRXL \reg_file_reg[9][15]  ( .D(n603), .CK(clk), .RN(n2276), .QN(n1825) );
  DFFRXL \reg_file_reg[9][14]  ( .D(n604), .CK(clk), .RN(n2277), .QN(n1824) );
  DFFRXL \reg_file_reg[9][13]  ( .D(n605), .CK(clk), .RN(n2277), .QN(n1823) );
  DFFRXL \reg_file_reg[9][12]  ( .D(n606), .CK(clk), .RN(n2278), .QN(n1822) );
  DFFRXL \reg_file_reg[9][11]  ( .D(n607), .CK(clk), .RN(n2278), .QN(n1821) );
  DFFRXL \reg_file_reg[9][10]  ( .D(n608), .CK(clk), .RN(n2279), .QN(n1820) );
  DFFRXL \reg_file_reg[9][9]  ( .D(n609), .CK(clk), .RN(n2279), .QN(n1819) );
  DFFRXL \reg_file_reg[9][8]  ( .D(n610), .CK(clk), .RN(n2280), .QN(n1818) );
  DFFRXL \reg_file_reg[9][7]  ( .D(n611), .CK(clk), .RN(n2280), .QN(n1817) );
  DFFRXL \reg_file_reg[9][6]  ( .D(n612), .CK(clk), .RN(n2281), .QN(n1816) );
  DFFRXL \reg_file_reg[9][5]  ( .D(n613), .CK(clk), .RN(n2285), .QN(n1815) );
  DFFRXL \reg_file_reg[9][4]  ( .D(n614), .CK(clk), .RN(n2285), .QN(n1814) );
  DFFRXL \reg_file_reg[9][3]  ( .D(n615), .CK(clk), .RN(n2285), .QN(n1813) );
  DFFRXL \reg_file_reg[9][2]  ( .D(n616), .CK(clk), .RN(n2282), .QN(n1812) );
  DFFRXL \reg_file_reg[9][1]  ( .D(n617), .CK(clk), .RN(n2285), .QN(n1811) );
  DFFRXL \reg_file_reg[9][0]  ( .D(n618), .CK(clk), .RN(n2285), .QN(n1810) );
  DFFRXL \reg_file_reg[10][31]  ( .D(n619), .CK(clk), .RN(n2274), .QN(n1809)
         );
  DFFRXL \reg_file_reg[10][30]  ( .D(n620), .CK(clk), .RN(n2277), .QN(n1808)
         );
  DFFRXL \reg_file_reg[10][29]  ( .D(n621), .CK(clk), .RN(n2271), .QN(n1807)
         );
  DFFRXL \reg_file_reg[10][28]  ( .D(n622), .CK(clk), .RN(n2271), .QN(n1806)
         );
  DFFRXL \reg_file_reg[10][27]  ( .D(n623), .CK(clk), .RN(n2272), .QN(n1805)
         );
  DFFRXL \reg_file_reg[10][26]  ( .D(n624), .CK(clk), .RN(n2273), .QN(n1804)
         );
  DFFRXL \reg_file_reg[10][25]  ( .D(n625), .CK(clk), .RN(n2273), .QN(n1803)
         );
  DFFRXL \reg_file_reg[10][24]  ( .D(n626), .CK(clk), .RN(n2271), .QN(n1802)
         );
  DFFRXL \reg_file_reg[10][23]  ( .D(n627), .CK(clk), .RN(n2274), .QN(n1801)
         );
  DFFRXL \reg_file_reg[10][22]  ( .D(n628), .CK(clk), .RN(n2274), .QN(n1800)
         );
  DFFRXL \reg_file_reg[10][21]  ( .D(n629), .CK(clk), .RN(n2274), .QN(n1799)
         );
  DFFRXL \reg_file_reg[10][20]  ( .D(n630), .CK(clk), .RN(n2274), .QN(n1798)
         );
  DFFRXL \reg_file_reg[10][19]  ( .D(n631), .CK(clk), .RN(n2277), .QN(n1797)
         );
  DFFRXL \reg_file_reg[10][18]  ( .D(n632), .CK(clk), .RN(n2285), .QN(n1796)
         );
  DFFRXL \reg_file_reg[10][17]  ( .D(n633), .CK(clk), .RN(n2275), .QN(n1795)
         );
  DFFRXL \reg_file_reg[10][16]  ( .D(n634), .CK(clk), .RN(n2275), .QN(n1794)
         );
  DFFRXL \reg_file_reg[10][15]  ( .D(n635), .CK(clk), .RN(n2276), .QN(n1793)
         );
  DFFRXL \reg_file_reg[10][14]  ( .D(n636), .CK(clk), .RN(n2277), .QN(n1792)
         );
  DFFRXL \reg_file_reg[10][13]  ( .D(n637), .CK(clk), .RN(n2277), .QN(n1791)
         );
  DFFRXL \reg_file_reg[10][12]  ( .D(n638), .CK(clk), .RN(n2278), .QN(n1790)
         );
  DFFRXL \reg_file_reg[10][11]  ( .D(n639), .CK(clk), .RN(n2278), .QN(n1789)
         );
  DFFRXL \reg_file_reg[10][10]  ( .D(n640), .CK(clk), .RN(n2279), .QN(n1788)
         );
  DFFRXL \reg_file_reg[10][9]  ( .D(n641), .CK(clk), .RN(n2279), .QN(n1787) );
  DFFRXL \reg_file_reg[10][8]  ( .D(n642), .CK(clk), .RN(n2280), .QN(n1786) );
  DFFRXL \reg_file_reg[10][7]  ( .D(n643), .CK(clk), .RN(n2280), .QN(n1785) );
  DFFRXL \reg_file_reg[10][6]  ( .D(n644), .CK(clk), .RN(n2281), .QN(n1784) );
  DFFRXL \reg_file_reg[10][5]  ( .D(n645), .CK(clk), .RN(n2285), .QN(n1783) );
  DFFRXL \reg_file_reg[10][4]  ( .D(n646), .CK(clk), .RN(n2285), .QN(n1782) );
  DFFRXL \reg_file_reg[10][3]  ( .D(n647), .CK(clk), .RN(n2285), .QN(n1781) );
  DFFRXL \reg_file_reg[10][2]  ( .D(n648), .CK(clk), .RN(n2281), .QN(n1780) );
  DFFRXL \reg_file_reg[10][1]  ( .D(n649), .CK(clk), .RN(n2285), .QN(n1779) );
  DFFRXL \reg_file_reg[10][0]  ( .D(n650), .CK(clk), .RN(n2285), .QN(n1778) );
  DFFRXL \reg_file_reg[11][31]  ( .D(n651), .CK(clk), .RN(n2273), .QN(n1777)
         );
  DFFRXL \reg_file_reg[11][30]  ( .D(n652), .CK(clk), .RN(n2272), .QN(n1776)
         );
  DFFRXL \reg_file_reg[11][29]  ( .D(n653), .CK(clk), .RN(n2271), .QN(n1775)
         );
  DFFRXL \reg_file_reg[11][28]  ( .D(n654), .CK(clk), .RN(n2271), .QN(n1774)
         );
  DFFRXL \reg_file_reg[11][27]  ( .D(n655), .CK(clk), .RN(n2272), .QN(n1773)
         );
  DFFRXL \reg_file_reg[11][26]  ( .D(n656), .CK(clk), .RN(n2273), .QN(n1772)
         );
  DFFRXL \reg_file_reg[11][25]  ( .D(n657), .CK(clk), .RN(n2273), .QN(n1771)
         );
  DFFRXL \reg_file_reg[11][24]  ( .D(n658), .CK(clk), .RN(n2277), .QN(n1770)
         );
  DFFRXL \reg_file_reg[11][23]  ( .D(n659), .CK(clk), .RN(n2273), .QN(n1769)
         );
  DFFRXL \reg_file_reg[11][22]  ( .D(n660), .CK(clk), .RN(n2274), .QN(n1768)
         );
  DFFRXL \reg_file_reg[11][21]  ( .D(n661), .CK(clk), .RN(n2274), .QN(n1767)
         );
  DFFRXL \reg_file_reg[11][20]  ( .D(n662), .CK(clk), .RN(n2273), .QN(n1766)
         );
  DFFRXL \reg_file_reg[11][19]  ( .D(n663), .CK(clk), .RN(n2272), .QN(n1765)
         );
  DFFRXL \reg_file_reg[11][18]  ( .D(n664), .CK(clk), .RN(n2285), .QN(n1764)
         );
  DFFRXL \reg_file_reg[11][17]  ( .D(n665), .CK(clk), .RN(n2275), .QN(n1763)
         );
  DFFRXL \reg_file_reg[11][16]  ( .D(n666), .CK(clk), .RN(n2275), .QN(n1762)
         );
  DFFRXL \reg_file_reg[11][15]  ( .D(n667), .CK(clk), .RN(n2276), .QN(n1761)
         );
  DFFRXL \reg_file_reg[11][14]  ( .D(n668), .CK(clk), .RN(n2277), .QN(n1760)
         );
  DFFRXL \reg_file_reg[11][13]  ( .D(n669), .CK(clk), .RN(n2277), .QN(n1759)
         );
  DFFRXL \reg_file_reg[11][12]  ( .D(n670), .CK(clk), .RN(n2278), .QN(n1758)
         );
  DFFRXL \reg_file_reg[11][11]  ( .D(n671), .CK(clk), .RN(n2278), .QN(n1757)
         );
  DFFRXL \reg_file_reg[11][10]  ( .D(n672), .CK(clk), .RN(n2279), .QN(n1756)
         );
  DFFRXL \reg_file_reg[11][9]  ( .D(n673), .CK(clk), .RN(n2279), .QN(n1755) );
  DFFRXL \reg_file_reg[11][8]  ( .D(n674), .CK(clk), .RN(n2280), .QN(n1754) );
  DFFRXL \reg_file_reg[11][7]  ( .D(n675), .CK(clk), .RN(n2280), .QN(n1753) );
  DFFRXL \reg_file_reg[11][6]  ( .D(n676), .CK(clk), .RN(n2281), .QN(n1752) );
  DFFRXL \reg_file_reg[11][5]  ( .D(n677), .CK(clk), .RN(n2285), .QN(n1751) );
  DFFRXL \reg_file_reg[11][4]  ( .D(n678), .CK(clk), .RN(n2285), .QN(n1750) );
  DFFRXL \reg_file_reg[11][3]  ( .D(n679), .CK(clk), .RN(n2285), .QN(n1749) );
  DFFRXL \reg_file_reg[11][2]  ( .D(n680), .CK(clk), .RN(n2281), .QN(n1748) );
  DFFRXL \reg_file_reg[11][1]  ( .D(n681), .CK(clk), .RN(n2285), .QN(n1747) );
  DFFRXL \reg_file_reg[11][0]  ( .D(n682), .CK(clk), .RN(n2285), .QN(n1746) );
  DFFRXL \reg_file_reg[12][31]  ( .D(n683), .CK(clk), .RN(n2276), .QN(n1745)
         );
  DFFRXL \reg_file_reg[12][30]  ( .D(n684), .CK(clk), .RN(n2277), .QN(n1744)
         );
  DFFRXL \reg_file_reg[12][29]  ( .D(n685), .CK(clk), .RN(n2271), .QN(n1743)
         );
  DFFRXL \reg_file_reg[12][28]  ( .D(n686), .CK(clk), .RN(n2271), .QN(n1742)
         );
  DFFRXL \reg_file_reg[12][27]  ( .D(n687), .CK(clk), .RN(n2272), .QN(n1741)
         );
  DFFRXL \reg_file_reg[12][26]  ( .D(n688), .CK(clk), .RN(n2273), .QN(n1740)
         );
  DFFRXL \reg_file_reg[12][25]  ( .D(n689), .CK(clk), .RN(n2273), .QN(n1739)
         );
  DFFRXL \reg_file_reg[12][24]  ( .D(n690), .CK(clk), .RN(n2272), .QN(n1738)
         );
  DFFRXL \reg_file_reg[12][23]  ( .D(n691), .CK(clk), .RN(n2276), .QN(n1737)
         );
  DFFRXL \reg_file_reg[12][22]  ( .D(n692), .CK(clk), .RN(n2274), .QN(n1736)
         );
  DFFRXL \reg_file_reg[12][21]  ( .D(n693), .CK(clk), .RN(n2274), .QN(n1735)
         );
  DFFRXL \reg_file_reg[12][20]  ( .D(n694), .CK(clk), .RN(n2281), .QN(n1734)
         );
  DFFRXL \reg_file_reg[12][19]  ( .D(n695), .CK(clk), .RN(n2276), .QN(n1733)
         );
  DFFRXL \reg_file_reg[12][18]  ( .D(n696), .CK(clk), .RN(n2285), .QN(n1732)
         );
  DFFRXL \reg_file_reg[12][17]  ( .D(n697), .CK(clk), .RN(n2275), .QN(n1731)
         );
  DFFRXL \reg_file_reg[12][16]  ( .D(n698), .CK(clk), .RN(n2275), .QN(n1730)
         );
  DFFRXL \reg_file_reg[12][15]  ( .D(n699), .CK(clk), .RN(n2276), .QN(n1729)
         );
  DFFRXL \reg_file_reg[12][14]  ( .D(n700), .CK(clk), .RN(n2277), .QN(n1728)
         );
  DFFRXL \reg_file_reg[12][13]  ( .D(n701), .CK(clk), .RN(n2277), .QN(n1727)
         );
  DFFRXL \reg_file_reg[12][12]  ( .D(n702), .CK(clk), .RN(n2278), .QN(n1726)
         );
  DFFRXL \reg_file_reg[12][11]  ( .D(n703), .CK(clk), .RN(n2278), .QN(n1725)
         );
  DFFRXL \reg_file_reg[12][10]  ( .D(n704), .CK(clk), .RN(n2279), .QN(n1724)
         );
  DFFRXL \reg_file_reg[12][9]  ( .D(n705), .CK(clk), .RN(n2279), .QN(n1723) );
  DFFRXL \reg_file_reg[12][8]  ( .D(n706), .CK(clk), .RN(n2280), .QN(n1722) );
  DFFRXL \reg_file_reg[12][7]  ( .D(n707), .CK(clk), .RN(n2280), .QN(n1721) );
  DFFRXL \reg_file_reg[12][6]  ( .D(n708), .CK(clk), .RN(n2281), .QN(n1720) );
  DFFRXL \reg_file_reg[12][5]  ( .D(n709), .CK(clk), .RN(n2285), .QN(n1719) );
  DFFRXL \reg_file_reg[12][4]  ( .D(n710), .CK(clk), .RN(n2285), .QN(n1718) );
  DFFRXL \reg_file_reg[12][3]  ( .D(n711), .CK(clk), .RN(n2285), .QN(n1717) );
  DFFRXL \reg_file_reg[12][2]  ( .D(n712), .CK(clk), .RN(n2281), .QN(n1716) );
  DFFRXL \reg_file_reg[12][1]  ( .D(n713), .CK(clk), .RN(n2285), .QN(n1715) );
  DFFRXL \reg_file_reg[12][0]  ( .D(n714), .CK(clk), .RN(n2285), .QN(n1714) );
  DFFRXL \reg_file_reg[13][31]  ( .D(n715), .CK(clk), .RN(n2275), .QN(n1713)
         );
  DFFRXL \reg_file_reg[13][30]  ( .D(n716), .CK(clk), .RN(n2280), .QN(n1712)
         );
  DFFRXL \reg_file_reg[13][29]  ( .D(n717), .CK(clk), .RN(n2271), .QN(n1711)
         );
  DFFRXL \reg_file_reg[13][28]  ( .D(n718), .CK(clk), .RN(n2271), .QN(n1710)
         );
  DFFRXL \reg_file_reg[13][27]  ( .D(n719), .CK(clk), .RN(n2272), .QN(n1709)
         );
  DFFRXL \reg_file_reg[13][26]  ( .D(n720), .CK(clk), .RN(n2272), .QN(n1708)
         );
  DFFRXL \reg_file_reg[13][25]  ( .D(n721), .CK(clk), .RN(n2273), .QN(n1707)
         );
  DFFRXL \reg_file_reg[13][24]  ( .D(n722), .CK(clk), .RN(n2276), .QN(n1706)
         );
  DFFRXL \reg_file_reg[13][23]  ( .D(n723), .CK(clk), .RN(n2275), .QN(n1705)
         );
  DFFRXL \reg_file_reg[13][22]  ( .D(n724), .CK(clk), .RN(n2274), .QN(n1704)
         );
  DFFRXL \reg_file_reg[13][21]  ( .D(n725), .CK(clk), .RN(n2274), .QN(n1703)
         );
  DFFRXL \reg_file_reg[13][20]  ( .D(n726), .CK(clk), .RN(n2275), .QN(n1702)
         );
  DFFRXL \reg_file_reg[13][19]  ( .D(n727), .CK(clk), .RN(n2280), .QN(n1701)
         );
  DFFRXL \reg_file_reg[13][18]  ( .D(n728), .CK(clk), .RN(n2285), .QN(n1700)
         );
  DFFRXL \reg_file_reg[13][17]  ( .D(n729), .CK(clk), .RN(n2275), .QN(n1699)
         );
  DFFRXL \reg_file_reg[13][16]  ( .D(n730), .CK(clk), .RN(n2275), .QN(n1698)
         );
  DFFRXL \reg_file_reg[13][15]  ( .D(n731), .CK(clk), .RN(n2276), .QN(n1697)
         );
  DFFRXL \reg_file_reg[13][14]  ( .D(n732), .CK(clk), .RN(n2277), .QN(n1696)
         );
  DFFRXL \reg_file_reg[13][13]  ( .D(n733), .CK(clk), .RN(n2277), .QN(n1695)
         );
  DFFRXL \reg_file_reg[13][12]  ( .D(n734), .CK(clk), .RN(n2278), .QN(n1694)
         );
  DFFRXL \reg_file_reg[13][11]  ( .D(n735), .CK(clk), .RN(n2278), .QN(n1693)
         );
  DFFRXL \reg_file_reg[13][10]  ( .D(n736), .CK(clk), .RN(n2279), .QN(n1692)
         );
  DFFRXL \reg_file_reg[13][9]  ( .D(n737), .CK(clk), .RN(n2279), .QN(n1691) );
  DFFRXL \reg_file_reg[13][8]  ( .D(n738), .CK(clk), .RN(n2280), .QN(n1690) );
  DFFRXL \reg_file_reg[13][7]  ( .D(n739), .CK(clk), .RN(n2280), .QN(n1689) );
  DFFRXL \reg_file_reg[13][6]  ( .D(n740), .CK(clk), .RN(n2281), .QN(n1688) );
  DFFRXL \reg_file_reg[13][5]  ( .D(n741), .CK(clk), .RN(n2285), .QN(n1687) );
  DFFRXL \reg_file_reg[13][4]  ( .D(n742), .CK(clk), .RN(n2285), .QN(n1686) );
  DFFRXL \reg_file_reg[13][3]  ( .D(n743), .CK(clk), .RN(n2284), .QN(n1685) );
  DFFRXL \reg_file_reg[13][2]  ( .D(n744), .CK(clk), .RN(n2281), .QN(n1684) );
  DFFRXL \reg_file_reg[13][1]  ( .D(n745), .CK(clk), .RN(n2284), .QN(n1683) );
  DFFRXL \reg_file_reg[13][0]  ( .D(n746), .CK(clk), .RN(n2284), .QN(n1682) );
  DFFRXL \reg_file_reg[14][31]  ( .D(n747), .CK(clk), .RN(n2281), .QN(n1681)
         );
  DFFRXL \reg_file_reg[14][30]  ( .D(n748), .CK(clk), .RN(n2283), .QN(n1680)
         );
  DFFRXL \reg_file_reg[14][29]  ( .D(n749), .CK(clk), .RN(n2271), .QN(n1679)
         );
  DFFRXL \reg_file_reg[14][28]  ( .D(n750), .CK(clk), .RN(n2271), .QN(n1678)
         );
  DFFRXL \reg_file_reg[14][27]  ( .D(n751), .CK(clk), .RN(n2272), .QN(n1677)
         );
  DFFRXL \reg_file_reg[14][26]  ( .D(n752), .CK(clk), .RN(n2272), .QN(n1676)
         );
  DFFRXL \reg_file_reg[14][25]  ( .D(n753), .CK(clk), .RN(n2273), .QN(n1675)
         );
  DFFRXL \reg_file_reg[14][24]  ( .D(n754), .CK(clk), .RN(n2280), .QN(n1674)
         );
  DFFRXL \reg_file_reg[14][23]  ( .D(n755), .CK(clk), .RN(n2281), .QN(n1673)
         );
  DFFRXL \reg_file_reg[14][22]  ( .D(n756), .CK(clk), .RN(n2274), .QN(n1672)
         );
  DFFRXL \reg_file_reg[14][21]  ( .D(n757), .CK(clk), .RN(n2274), .QN(n1671)
         );
  DFFRXL \reg_file_reg[14][20]  ( .D(n758), .CK(clk), .RN(n2283), .QN(n1670)
         );
  DFFRXL \reg_file_reg[14][19]  ( .D(n759), .CK(clk), .RN(n2284), .QN(n1669)
         );
  DFFRXL \reg_file_reg[14][18]  ( .D(n760), .CK(clk), .RN(n2284), .QN(n1668)
         );
  DFFRXL \reg_file_reg[14][17]  ( .D(n761), .CK(clk), .RN(n2275), .QN(n1667)
         );
  DFFRXL \reg_file_reg[14][16]  ( .D(n762), .CK(clk), .RN(n2275), .QN(n1666)
         );
  DFFRXL \reg_file_reg[14][15]  ( .D(n763), .CK(clk), .RN(n2276), .QN(n1665)
         );
  DFFRXL \reg_file_reg[14][14]  ( .D(n764), .CK(clk), .RN(n2277), .QN(n1664)
         );
  DFFRXL \reg_file_reg[14][13]  ( .D(n765), .CK(clk), .RN(n2277), .QN(n1663)
         );
  DFFRXL \reg_file_reg[14][12]  ( .D(n766), .CK(clk), .RN(n2278), .QN(n1662)
         );
  DFFRXL \reg_file_reg[14][11]  ( .D(n767), .CK(clk), .RN(n2278), .QN(n1661)
         );
  DFFRXL \reg_file_reg[14][10]  ( .D(n768), .CK(clk), .RN(n2279), .QN(n1660)
         );
  DFFRXL \reg_file_reg[14][9]  ( .D(n769), .CK(clk), .RN(n2279), .QN(n1659) );
  DFFRXL \reg_file_reg[14][8]  ( .D(n770), .CK(clk), .RN(n2280), .QN(n1658) );
  DFFRXL \reg_file_reg[14][7]  ( .D(n771), .CK(clk), .RN(n2280), .QN(n1657) );
  DFFRXL \reg_file_reg[14][6]  ( .D(n772), .CK(clk), .RN(n2281), .QN(n1656) );
  DFFRXL \reg_file_reg[14][5]  ( .D(n773), .CK(clk), .RN(n2284), .QN(n1655) );
  DFFRXL \reg_file_reg[14][4]  ( .D(n774), .CK(clk), .RN(n2284), .QN(n1654) );
  DFFRXL \reg_file_reg[14][3]  ( .D(n775), .CK(clk), .RN(n2284), .QN(n1653) );
  DFFRXL \reg_file_reg[14][2]  ( .D(n776), .CK(clk), .RN(n2281), .QN(n1652) );
  DFFRXL \reg_file_reg[14][1]  ( .D(n777), .CK(clk), .RN(n2284), .QN(n1651) );
  DFFRXL \reg_file_reg[14][0]  ( .D(n778), .CK(clk), .RN(n2284), .QN(n1650) );
  DFFRXL \reg_file_reg[15][31]  ( .D(n779), .CK(clk), .RN(n2283), .QN(n1649)
         );
  DFFRXL \reg_file_reg[15][30]  ( .D(n780), .CK(clk), .RN(n2284), .QN(n1648)
         );
  DFFRXL \reg_file_reg[15][29]  ( .D(n781), .CK(clk), .RN(n2271), .QN(n1647)
         );
  DFFRXL \reg_file_reg[15][28]  ( .D(n782), .CK(clk), .RN(n2271), .QN(n1646)
         );
  DFFRXL \reg_file_reg[15][27]  ( .D(n783), .CK(clk), .RN(n2272), .QN(n1645)
         );
  DFFRXL \reg_file_reg[15][26]  ( .D(n784), .CK(clk), .RN(n2272), .QN(n1644)
         );
  DFFRXL \reg_file_reg[15][25]  ( .D(n785), .CK(clk), .RN(n2273), .QN(n1643)
         );
  DFFRXL \reg_file_reg[15][24]  ( .D(n786), .CK(clk), .RN(n2283), .QN(n1642)
         );
  DFFRXL \reg_file_reg[15][23]  ( .D(n787), .CK(clk), .RN(n2284), .QN(n1641)
         );
  DFFRXL \reg_file_reg[15][22]  ( .D(n788), .CK(clk), .RN(n2274), .QN(n1640)
         );
  DFFRXL \reg_file_reg[15][21]  ( .D(n789), .CK(clk), .RN(n2274), .QN(n1639)
         );
  DFFRXL \reg_file_reg[15][20]  ( .D(n790), .CK(clk), .RN(n2282), .QN(n1638)
         );
  DFFRXL \reg_file_reg[15][19]  ( .D(n791), .CK(clk), .RN(n2278), .QN(n1637)
         );
  DFFRXL \reg_file_reg[15][18]  ( .D(n792), .CK(clk), .RN(n2284), .QN(n1636)
         );
  DFFRXL \reg_file_reg[15][17]  ( .D(n793), .CK(clk), .RN(n2275), .QN(n1635)
         );
  DFFRXL \reg_file_reg[15][16]  ( .D(n794), .CK(clk), .RN(n2275), .QN(n1634)
         );
  DFFRXL \reg_file_reg[15][15]  ( .D(n795), .CK(clk), .RN(n2276), .QN(n1633)
         );
  DFFRXL \reg_file_reg[15][14]  ( .D(n796), .CK(clk), .RN(n2277), .QN(n1632)
         );
  DFFRXL \reg_file_reg[15][13]  ( .D(n797), .CK(clk), .RN(n2277), .QN(n1631)
         );
  DFFRXL \reg_file_reg[15][12]  ( .D(n798), .CK(clk), .RN(n2278), .QN(n1630)
         );
  DFFRXL \reg_file_reg[15][11]  ( .D(n799), .CK(clk), .RN(n2278), .QN(n1629)
         );
  DFFRXL \reg_file_reg[15][10]  ( .D(n800), .CK(clk), .RN(n2279), .QN(n1628)
         );
  DFFRXL \reg_file_reg[15][9]  ( .D(n801), .CK(clk), .RN(n2279), .QN(n1627) );
  DFFRXL \reg_file_reg[15][8]  ( .D(n802), .CK(clk), .RN(n2280), .QN(n1626) );
  DFFRXL \reg_file_reg[15][7]  ( .D(n803), .CK(clk), .RN(n2280), .QN(n1625) );
  DFFRXL \reg_file_reg[15][6]  ( .D(n804), .CK(clk), .RN(n2281), .QN(n1624) );
  DFFRXL \reg_file_reg[15][5]  ( .D(n805), .CK(clk), .RN(n2284), .QN(n1623) );
  DFFRXL \reg_file_reg[15][4]  ( .D(n806), .CK(clk), .RN(n2284), .QN(n1622) );
  DFFRXL \reg_file_reg[15][3]  ( .D(n807), .CK(clk), .RN(n2284), .QN(n1621) );
  DFFRXL \reg_file_reg[15][2]  ( .D(n808), .CK(clk), .RN(n2281), .QN(n1620) );
  DFFRXL \reg_file_reg[15][1]  ( .D(n809), .CK(clk), .RN(n2284), .QN(n1619) );
  DFFRXL \reg_file_reg[15][0]  ( .D(n810), .CK(clk), .RN(n2284), .QN(n1618) );
  DFFRXL \reg_file_reg[16][31]  ( .D(n811), .CK(clk), .RN(n2278), .QN(n1617)
         );
  DFFRXL \reg_file_reg[16][30]  ( .D(n812), .CK(clk), .RN(n2282), .QN(n1616)
         );
  DFFRXL \reg_file_reg[16][29]  ( .D(n813), .CK(clk), .RN(n2271), .QN(n1615)
         );
  DFFRXL \reg_file_reg[16][28]  ( .D(n814), .CK(clk), .RN(n2271), .QN(n1614)
         );
  DFFRXL \reg_file_reg[16][27]  ( .D(n815), .CK(clk), .RN(n2272), .QN(n1613)
         );
  DFFRXL \reg_file_reg[16][26]  ( .D(n816), .CK(clk), .RN(n2272), .QN(n1612)
         );
  DFFRXL \reg_file_reg[16][25]  ( .D(n817), .CK(clk), .RN(n2273), .QN(n1611)
         );
  DFFRXL \reg_file_reg[16][24]  ( .D(n818), .CK(clk), .RN(n2282), .QN(n1610)
         );
  DFFRXL \reg_file_reg[16][23]  ( .D(n819), .CK(clk), .RN(n2278), .QN(n1609)
         );
  DFFRXL \reg_file_reg[16][22]  ( .D(n820), .CK(clk), .RN(n2274), .QN(n1608)
         );
  DFFRXL \reg_file_reg[16][21]  ( .D(n821), .CK(clk), .RN(n2274), .QN(n1607)
         );
  DFFRXL \reg_file_reg[16][20]  ( .D(n822), .CK(clk), .RN(n2279), .QN(n1606)
         );
  DFFRXL \reg_file_reg[16][19]  ( .D(n823), .CK(clk), .RN(n2271), .QN(n1605)
         );
  DFFRXL \reg_file_reg[16][18]  ( .D(n824), .CK(clk), .RN(n2282), .QN(n1604)
         );
  DFFRXL \reg_file_reg[16][17]  ( .D(n825), .CK(clk), .RN(n2275), .QN(n1603)
         );
  DFFRXL \reg_file_reg[16][16]  ( .D(n826), .CK(clk), .RN(n2275), .QN(n1602)
         );
  DFFRXL \reg_file_reg[16][15]  ( .D(n827), .CK(clk), .RN(n2276), .QN(n1601)
         );
  DFFRXL \reg_file_reg[16][14]  ( .D(n828), .CK(clk), .RN(n2276), .QN(n1600)
         );
  DFFRXL \reg_file_reg[16][13]  ( .D(n829), .CK(clk), .RN(n2277), .QN(n1599)
         );
  DFFRXL \reg_file_reg[16][12]  ( .D(n830), .CK(clk), .RN(n2278), .QN(n1598)
         );
  DFFRXL \reg_file_reg[16][11]  ( .D(n831), .CK(clk), .RN(n2278), .QN(n1597)
         );
  DFFRXL \reg_file_reg[16][10]  ( .D(n832), .CK(clk), .RN(n2279), .QN(n1596)
         );
  DFFRXL \reg_file_reg[16][9]  ( .D(n833), .CK(clk), .RN(n2279), .QN(n1595) );
  DFFRXL \reg_file_reg[16][8]  ( .D(n834), .CK(clk), .RN(n2280), .QN(n1594) );
  DFFRXL \reg_file_reg[16][7]  ( .D(n835), .CK(clk), .RN(n2280), .QN(n1593) );
  DFFRXL \reg_file_reg[16][6]  ( .D(n836), .CK(clk), .RN(n2281), .QN(n1592) );
  DFFRXL \reg_file_reg[16][5]  ( .D(n837), .CK(clk), .RN(n2282), .QN(n1591) );
  DFFRXL \reg_file_reg[16][4]  ( .D(n838), .CK(clk), .RN(n2282), .QN(n1590) );
  DFFRXL \reg_file_reg[16][3]  ( .D(n839), .CK(clk), .RN(n2282), .QN(n1589) );
  DFFRXL \reg_file_reg[16][2]  ( .D(n840), .CK(clk), .RN(n2281), .QN(n1588) );
  DFFRXL \reg_file_reg[16][1]  ( .D(n841), .CK(clk), .RN(n2282), .QN(n1587) );
  DFFRXL \reg_file_reg[16][0]  ( .D(n842), .CK(clk), .RN(n2282), .QN(n1586) );
  DFFRXL \reg_file_reg[17][31]  ( .D(n843), .CK(clk), .RN(n2279), .QN(n1585)
         );
  DFFRXL \reg_file_reg[17][30]  ( .D(n844), .CK(clk), .RN(n2271), .QN(n1584)
         );
  DFFRXL \reg_file_reg[17][29]  ( .D(n845), .CK(clk), .RN(n2271), .QN(n1583)
         );
  DFFRXL \reg_file_reg[17][28]  ( .D(n846), .CK(clk), .RN(n2271), .QN(n1582)
         );
  DFFRXL \reg_file_reg[17][27]  ( .D(n847), .CK(clk), .RN(n2272), .QN(n1581)
         );
  DFFRXL \reg_file_reg[17][26]  ( .D(n848), .CK(clk), .RN(n2272), .QN(n1580)
         );
  DFFRXL \reg_file_reg[17][25]  ( .D(n849), .CK(clk), .RN(n2273), .QN(n1579)
         );
  DFFRXL \reg_file_reg[17][24]  ( .D(n850), .CK(clk), .RN(n2279), .QN(n1578)
         );
  DFFRXL \reg_file_reg[17][23]  ( .D(n851), .CK(clk), .RN(n2271), .QN(n1577)
         );
  DFFRXL \reg_file_reg[17][22]  ( .D(n852), .CK(clk), .RN(n2274), .QN(n1576)
         );
  DFFRXL \reg_file_reg[17][21]  ( .D(n853), .CK(clk), .RN(n2274), .QN(n1575)
         );
  DFFRXL \reg_file_reg[17][20]  ( .D(n854), .CK(clk), .RN(n2274), .QN(n1574)
         );
  DFFRXL \reg_file_reg[17][19]  ( .D(n855), .CK(clk), .RN(n2277), .QN(n1573)
         );
  DFFRXL \reg_file_reg[17][18]  ( .D(n856), .CK(clk), .RN(n2282), .QN(n1572)
         );
  DFFRXL \reg_file_reg[17][17]  ( .D(n857), .CK(clk), .RN(n2275), .QN(n1571)
         );
  DFFRXL \reg_file_reg[17][16]  ( .D(n858), .CK(clk), .RN(n2275), .QN(n1570)
         );
  DFFRXL \reg_file_reg[17][15]  ( .D(n859), .CK(clk), .RN(n2276), .QN(n1569)
         );
  DFFRXL \reg_file_reg[17][14]  ( .D(n860), .CK(clk), .RN(n2276), .QN(n1568)
         );
  DFFRXL \reg_file_reg[17][13]  ( .D(n861), .CK(clk), .RN(n2277), .QN(n1567)
         );
  DFFRXL \reg_file_reg[17][12]  ( .D(n862), .CK(clk), .RN(n2278), .QN(n1566)
         );
  DFFRXL \reg_file_reg[17][11]  ( .D(n863), .CK(clk), .RN(n2278), .QN(n1565)
         );
  DFFRXL \reg_file_reg[17][10]  ( .D(n864), .CK(clk), .RN(n2279), .QN(n1564)
         );
  DFFRXL \reg_file_reg[17][9]  ( .D(n865), .CK(clk), .RN(n2279), .QN(n1563) );
  DFFRXL \reg_file_reg[17][8]  ( .D(n866), .CK(clk), .RN(n2280), .QN(n1562) );
  DFFRXL \reg_file_reg[17][7]  ( .D(n867), .CK(clk), .RN(n2280), .QN(n1561) );
  DFFRXL \reg_file_reg[17][6]  ( .D(n868), .CK(clk), .RN(n2281), .QN(n1560) );
  DFFRXL \reg_file_reg[17][5]  ( .D(n869), .CK(clk), .RN(n2282), .QN(n1559) );
  DFFRXL \reg_file_reg[17][4]  ( .D(n870), .CK(clk), .RN(n2282), .QN(n1558) );
  DFFRXL \reg_file_reg[17][3]  ( .D(n871), .CK(clk), .RN(n2282), .QN(n1557) );
  DFFRXL \reg_file_reg[17][2]  ( .D(n872), .CK(clk), .RN(n2281), .QN(n1556) );
  DFFRXL \reg_file_reg[17][1]  ( .D(n873), .CK(clk), .RN(n2282), .QN(n1555) );
  DFFRXL \reg_file_reg[17][0]  ( .D(n874), .CK(clk), .RN(n2282), .QN(n1554) );
  DFFRXL \reg_file_reg[18][31]  ( .D(n875), .CK(clk), .RN(n2274), .QN(n1553)
         );
  DFFRXL \reg_file_reg[18][30]  ( .D(n876), .CK(clk), .RN(n2277), .QN(n1552)
         );
  DFFRXL \reg_file_reg[18][29]  ( .D(n877), .CK(clk), .RN(n2271), .QN(n1551)
         );
  DFFRXL \reg_file_reg[18][28]  ( .D(n878), .CK(clk), .RN(n2271), .QN(n1550)
         );
  DFFRXL \reg_file_reg[18][27]  ( .D(n879), .CK(clk), .RN(n2272), .QN(n1549)
         );
  DFFRXL \reg_file_reg[18][26]  ( .D(n880), .CK(clk), .RN(n2272), .QN(n1548)
         );
  DFFRXL \reg_file_reg[18][25]  ( .D(n881), .CK(clk), .RN(n2273), .QN(n1547)
         );
  DFFRXL \reg_file_reg[18][24]  ( .D(n882), .CK(clk), .RN(n2274), .QN(n1546)
         );
  DFFRXL \reg_file_reg[18][23]  ( .D(n883), .CK(clk), .RN(n2277), .QN(n1545)
         );
  DFFRXL \reg_file_reg[18][22]  ( .D(n884), .CK(clk), .RN(n2274), .QN(n1544)
         );
  DFFRXL \reg_file_reg[18][21]  ( .D(n885), .CK(clk), .RN(n2274), .QN(n1543)
         );
  DFFRXL \reg_file_reg[18][20]  ( .D(n886), .CK(clk), .RN(n2273), .QN(n1542)
         );
  DFFRXL \reg_file_reg[18][19]  ( .D(n887), .CK(clk), .RN(n2272), .QN(n1541)
         );
  DFFRXL \reg_file_reg[18][18]  ( .D(n888), .CK(clk), .RN(n2282), .QN(n1540)
         );
  DFFRXL \reg_file_reg[18][17]  ( .D(n889), .CK(clk), .RN(n2275), .QN(n1539)
         );
  DFFRXL \reg_file_reg[18][16]  ( .D(n890), .CK(clk), .RN(n2275), .QN(n1538)
         );
  DFFRXL \reg_file_reg[18][15]  ( .D(n891), .CK(clk), .RN(n2276), .QN(n1537)
         );
  DFFRXL \reg_file_reg[18][14]  ( .D(n892), .CK(clk), .RN(n2276), .QN(n1536)
         );
  DFFRXL \reg_file_reg[18][13]  ( .D(n893), .CK(clk), .RN(n2277), .QN(n1535)
         );
  DFFRXL \reg_file_reg[18][12]  ( .D(n894), .CK(clk), .RN(n2278), .QN(n1534)
         );
  DFFRXL \reg_file_reg[18][11]  ( .D(n895), .CK(clk), .RN(n2278), .QN(n1533)
         );
  DFFRXL \reg_file_reg[18][10]  ( .D(n896), .CK(clk), .RN(n2279), .QN(n1532)
         );
  DFFRXL \reg_file_reg[18][9]  ( .D(n897), .CK(clk), .RN(n2279), .QN(n1531) );
  DFFRXL \reg_file_reg[18][8]  ( .D(n898), .CK(clk), .RN(n2280), .QN(n1530) );
  DFFRXL \reg_file_reg[18][7]  ( .D(n899), .CK(clk), .RN(n2280), .QN(n1529) );
  DFFRXL \reg_file_reg[18][6]  ( .D(n900), .CK(clk), .RN(n2281), .QN(n1528) );
  DFFRXL \reg_file_reg[18][5]  ( .D(n901), .CK(clk), .RN(n2282), .QN(n1527) );
  DFFRXL \reg_file_reg[18][4]  ( .D(n902), .CK(clk), .RN(n2282), .QN(n1526) );
  DFFRXL \reg_file_reg[18][3]  ( .D(n903), .CK(clk), .RN(n2282), .QN(n1525) );
  DFFRXL \reg_file_reg[18][2]  ( .D(n904), .CK(clk), .RN(n2281), .QN(n1524) );
  DFFRXL \reg_file_reg[18][1]  ( .D(n905), .CK(clk), .RN(n2282), .QN(n1523) );
  DFFRXL \reg_file_reg[18][0]  ( .D(n906), .CK(clk), .RN(n2282), .QN(n1522) );
  DFFRXL \reg_file_reg[19][31]  ( .D(n907), .CK(clk), .RN(n2273), .QN(n1521)
         );
  DFFRXL \reg_file_reg[19][30]  ( .D(n908), .CK(clk), .RN(n2272), .QN(n1520)
         );
  DFFRXL \reg_file_reg[19][29]  ( .D(n909), .CK(clk), .RN(n2271), .QN(n1519)
         );
  DFFRXL \reg_file_reg[19][28]  ( .D(n910), .CK(clk), .RN(n2271), .QN(n1518)
         );
  DFFRXL \reg_file_reg[19][27]  ( .D(n911), .CK(clk), .RN(n2272), .QN(n1517)
         );
  DFFRXL \reg_file_reg[19][26]  ( .D(n912), .CK(clk), .RN(n2272), .QN(n1516)
         );
  DFFRXL \reg_file_reg[19][25]  ( .D(n913), .CK(clk), .RN(n2273), .QN(n1515)
         );
  DFFRXL \reg_file_reg[19][24]  ( .D(n914), .CK(clk), .RN(n2273), .QN(n1514)
         );
  DFFRXL \reg_file_reg[19][23]  ( .D(n915), .CK(clk), .RN(n2273), .QN(n1513)
         );
  DFFRXL \reg_file_reg[19][22]  ( .D(n916), .CK(clk), .RN(n2274), .QN(n1512)
         );
  DFFRXL \reg_file_reg[19][21]  ( .D(n917), .CK(clk), .RN(n2274), .QN(n1511)
         );
  DFFRXL \reg_file_reg[19][20]  ( .D(n918), .CK(clk), .RN(n2281), .QN(n1510)
         );
  DFFRXL \reg_file_reg[19][19]  ( .D(n919), .CK(clk), .RN(n2276), .QN(n1509)
         );
  DFFRXL \reg_file_reg[19][18]  ( .D(n920), .CK(clk), .RN(n2282), .QN(n1508)
         );
  DFFRXL \reg_file_reg[19][17]  ( .D(n921), .CK(clk), .RN(n2275), .QN(n1507)
         );
  DFFRXL \reg_file_reg[19][16]  ( .D(n922), .CK(clk), .RN(n2275), .QN(n1506)
         );
  DFFRXL \reg_file_reg[19][15]  ( .D(n923), .CK(clk), .RN(n2276), .QN(n1505)
         );
  DFFRXL \reg_file_reg[19][14]  ( .D(n924), .CK(clk), .RN(n2276), .QN(n1504)
         );
  DFFRXL \reg_file_reg[19][13]  ( .D(n925), .CK(clk), .RN(n2277), .QN(n1503)
         );
  DFFRXL \reg_file_reg[19][12]  ( .D(n926), .CK(clk), .RN(n2278), .QN(n1502)
         );
  DFFRXL \reg_file_reg[19][11]  ( .D(n927), .CK(clk), .RN(n2278), .QN(n1501)
         );
  DFFRXL \reg_file_reg[19][10]  ( .D(n928), .CK(clk), .RN(n2279), .QN(n1500)
         );
  DFFRXL \reg_file_reg[19][9]  ( .D(n929), .CK(clk), .RN(n2279), .QN(n1499) );
  DFFRXL \reg_file_reg[19][8]  ( .D(n930), .CK(clk), .RN(n2280), .QN(n1498) );
  DFFRXL \reg_file_reg[19][7]  ( .D(n931), .CK(clk), .RN(n2280), .QN(n1497) );
  DFFRXL \reg_file_reg[19][6]  ( .D(n932), .CK(clk), .RN(n2281), .QN(n1496) );
  DFFRXL \reg_file_reg[19][5]  ( .D(n933), .CK(clk), .RN(n2282), .QN(n1495) );
  DFFRXL \reg_file_reg[19][4]  ( .D(n934), .CK(clk), .RN(n2282), .QN(n1494) );
  DFFRXL \reg_file_reg[19][3]  ( .D(n935), .CK(clk), .RN(n2282), .QN(n1493) );
  DFFRXL \reg_file_reg[19][2]  ( .D(n936), .CK(clk), .RN(n2281), .QN(n1492) );
  DFFRXL \reg_file_reg[19][1]  ( .D(n937), .CK(clk), .RN(n2282), .QN(n1491) );
  DFFRXL \reg_file_reg[19][0]  ( .D(n938), .CK(clk), .RN(n2282), .QN(n1490) );
  DFFRXL \reg_file_reg[20][31]  ( .D(n939), .CK(clk), .RN(n2276), .QN(n1489)
         );
  DFFRXL \reg_file_reg[20][30]  ( .D(n940), .CK(clk), .RN(n2273), .QN(n1488)
         );
  DFFRXL \reg_file_reg[20][29]  ( .D(n941), .CK(clk), .RN(n2271), .QN(n1487)
         );
  DFFRXL \reg_file_reg[20][28]  ( .D(n942), .CK(clk), .RN(n2271), .QN(n1486)
         );
  DFFRXL \reg_file_reg[20][27]  ( .D(n943), .CK(clk), .RN(n2272), .QN(n1485)
         );
  DFFRXL \reg_file_reg[20][26]  ( .D(n944), .CK(clk), .RN(n2272), .QN(n1484)
         );
  DFFRXL \reg_file_reg[20][25]  ( .D(n945), .CK(clk), .RN(n2273), .QN(n1483)
         );
  DFFRXL \reg_file_reg[20][24]  ( .D(n946), .CK(clk), .RN(n2273), .QN(n1482)
         );
  DFFRXL \reg_file_reg[20][23]  ( .D(n947), .CK(clk), .RN(n2272), .QN(n1481)
         );
  DFFRXL \reg_file_reg[20][22]  ( .D(n948), .CK(clk), .RN(n2274), .QN(n1480)
         );
  DFFRXL \reg_file_reg[20][21]  ( .D(n949), .CK(clk), .RN(n2274), .QN(n1479)
         );
  DFFRXL \reg_file_reg[20][20]  ( .D(n950), .CK(clk), .RN(n2275), .QN(n1478)
         );
  DFFRXL \reg_file_reg[20][19]  ( .D(n951), .CK(clk), .RN(n2280), .QN(n1477)
         );
  DFFRXL \reg_file_reg[20][18]  ( .D(n952), .CK(clk), .RN(n2282), .QN(n1476)
         );
  DFFRXL \reg_file_reg[20][17]  ( .D(n953), .CK(clk), .RN(n2275), .QN(n1475)
         );
  DFFRXL \reg_file_reg[20][16]  ( .D(n954), .CK(clk), .RN(n2275), .QN(n1474)
         );
  DFFRXL \reg_file_reg[20][15]  ( .D(n955), .CK(clk), .RN(n2276), .QN(n1473)
         );
  DFFRXL \reg_file_reg[20][14]  ( .D(n956), .CK(clk), .RN(n2276), .QN(n1472)
         );
  DFFRXL \reg_file_reg[20][13]  ( .D(n957), .CK(clk), .RN(n2277), .QN(n1471)
         );
  DFFRXL \reg_file_reg[20][12]  ( .D(n958), .CK(clk), .RN(n2278), .QN(n1470)
         );
  DFFRXL \reg_file_reg[20][11]  ( .D(n959), .CK(clk), .RN(n2278), .QN(n1469)
         );
  DFFRXL \reg_file_reg[20][10]  ( .D(n960), .CK(clk), .RN(n2279), .QN(n1468)
         );
  DFFRXL \reg_file_reg[20][9]  ( .D(n961), .CK(clk), .RN(n2279), .QN(n1467) );
  DFFRXL \reg_file_reg[20][8]  ( .D(n962), .CK(clk), .RN(n2280), .QN(n1466) );
  DFFRXL \reg_file_reg[20][7]  ( .D(n963), .CK(clk), .RN(n2280), .QN(n1465) );
  DFFRXL \reg_file_reg[20][6]  ( .D(n964), .CK(clk), .RN(n2281), .QN(n1464) );
  DFFRXL \reg_file_reg[20][5]  ( .D(n965), .CK(clk), .RN(n2282), .QN(n1463) );
  DFFRXL \reg_file_reg[20][4]  ( .D(n966), .CK(clk), .RN(n2282), .QN(n1462) );
  DFFRXL \reg_file_reg[20][3]  ( .D(n967), .CK(clk), .RN(n2282), .QN(n1461) );
  DFFRXL \reg_file_reg[20][2]  ( .D(n968), .CK(clk), .RN(n2281), .QN(n1460) );
  DFFRXL \reg_file_reg[20][1]  ( .D(n969), .CK(clk), .RN(n2282), .QN(n1459) );
  DFFRXL \reg_file_reg[20][0]  ( .D(n970), .CK(clk), .RN(n2282), .QN(n1458) );
  DFFRXL \reg_file_reg[21][31]  ( .D(n971), .CK(clk), .RN(n2275), .QN(n1457)
         );
  DFFRXL \reg_file_reg[21][30]  ( .D(n972), .CK(clk), .RN(n2280), .QN(n1456)
         );
  DFFRXL \reg_file_reg[21][29]  ( .D(n973), .CK(clk), .RN(n2271), .QN(n1455)
         );
  DFFRXL \reg_file_reg[21][28]  ( .D(n974), .CK(clk), .RN(n2271), .QN(n1454)
         );
  DFFRXL \reg_file_reg[21][27]  ( .D(n975), .CK(clk), .RN(n2272), .QN(n1453)
         );
  DFFRXL \reg_file_reg[21][26]  ( .D(n976), .CK(clk), .RN(n2272), .QN(n1452)
         );
  DFFRXL \reg_file_reg[21][25]  ( .D(n977), .CK(clk), .RN(n2273), .QN(n1451)
         );
  DFFRXL \reg_file_reg[21][24]  ( .D(n978), .CK(clk), .RN(n2273), .QN(n1450)
         );
  DFFRXL \reg_file_reg[21][23]  ( .D(n979), .CK(clk), .RN(n2276), .QN(n1449)
         );
  DFFRXL \reg_file_reg[21][22]  ( .D(n980), .CK(clk), .RN(n2274), .QN(n1448)
         );
  DFFRXL \reg_file_reg[21][21]  ( .D(n981), .CK(clk), .RN(n2274), .QN(n1447)
         );
  DFFRXL \reg_file_reg[21][20]  ( .D(n982), .CK(clk), .RN(n2283), .QN(n1446)
         );
  DFFRXL \reg_file_reg[21][19]  ( .D(n983), .CK(clk), .RN(n2284), .QN(n1445)
         );
  DFFRXL \reg_file_reg[21][18]  ( .D(n984), .CK(clk), .RN(n2283), .QN(n1444)
         );
  DFFRXL \reg_file_reg[21][17]  ( .D(n985), .CK(clk), .RN(n2275), .QN(n1443)
         );
  DFFRXL \reg_file_reg[21][16]  ( .D(n986), .CK(clk), .RN(n2275), .QN(n1442)
         );
  DFFRXL \reg_file_reg[21][15]  ( .D(n987), .CK(clk), .RN(n2276), .QN(n1441)
         );
  DFFRXL \reg_file_reg[21][14]  ( .D(n988), .CK(clk), .RN(n2276), .QN(n1440)
         );
  DFFRXL \reg_file_reg[21][13]  ( .D(n989), .CK(clk), .RN(n2277), .QN(n1439)
         );
  DFFRXL \reg_file_reg[21][12]  ( .D(n990), .CK(clk), .RN(n2278), .QN(n1438)
         );
  DFFRXL \reg_file_reg[21][11]  ( .D(n991), .CK(clk), .RN(n2278), .QN(n1437)
         );
  DFFRXL \reg_file_reg[21][10]  ( .D(n992), .CK(clk), .RN(n2279), .QN(n1436)
         );
  DFFRXL \reg_file_reg[21][9]  ( .D(n993), .CK(clk), .RN(n2279), .QN(n1435) );
  DFFRXL \reg_file_reg[21][8]  ( .D(n994), .CK(clk), .RN(n2280), .QN(n1434) );
  DFFRXL \reg_file_reg[21][7]  ( .D(n995), .CK(clk), .RN(n2280), .QN(n1433) );
  DFFRXL \reg_file_reg[21][6]  ( .D(n996), .CK(clk), .RN(n2281), .QN(n1432) );
  DFFRXL \reg_file_reg[21][5]  ( .D(n997), .CK(clk), .RN(n2283), .QN(n1431) );
  DFFRXL \reg_file_reg[21][4]  ( .D(n998), .CK(clk), .RN(n2283), .QN(n1430) );
  DFFRXL \reg_file_reg[21][3]  ( .D(n999), .CK(clk), .RN(n2283), .QN(n1429) );
  DFFRXL \reg_file_reg[21][2]  ( .D(n1000), .CK(clk), .RN(n2282), .QN(n1428)
         );
  DFFRXL \reg_file_reg[21][1]  ( .D(n1001), .CK(clk), .RN(n2283), .QN(n1427)
         );
  DFFRXL \reg_file_reg[21][0]  ( .D(n1002), .CK(clk), .RN(n2283), .QN(n1426)
         );
  DFFRXL \reg_file_reg[22][31]  ( .D(n1003), .CK(clk), .RN(n2281), .QN(n1425)
         );
  DFFRXL \reg_file_reg[22][30]  ( .D(n1004), .CK(clk), .RN(n2271), .QN(n1424)
         );
  DFFRXL \reg_file_reg[22][29]  ( .D(n1005), .CK(clk), .RN(n2271), .QN(n1423)
         );
  DFFRXL \reg_file_reg[22][28]  ( .D(n1006), .CK(clk), .RN(n2272), .QN(n1422)
         );
  DFFRXL \reg_file_reg[22][27]  ( .D(n1007), .CK(clk), .RN(n2272), .QN(n1421)
         );
  DFFRXL \reg_file_reg[22][26]  ( .D(n1008), .CK(clk), .RN(n2273), .QN(n1420)
         );
  DFFRXL \reg_file_reg[22][25]  ( .D(n1009), .CK(clk), .RN(n2273), .QN(n1419)
         );
  DFFRXL \reg_file_reg[22][24]  ( .D(n1010), .CK(clk), .RN(n2275), .QN(n1418)
         );
  DFFRXL \reg_file_reg[22][23]  ( .D(n1011), .CK(clk), .RN(n2274), .QN(n1417)
         );
  DFFRXL \reg_file_reg[22][22]  ( .D(n1012), .CK(clk), .RN(n2274), .QN(n1416)
         );
  DFFRXL \reg_file_reg[22][21]  ( .D(n1013), .CK(clk), .RN(n2282), .QN(n1415)
         );
  DFFRXL \reg_file_reg[22][20]  ( .D(n1014), .CK(clk), .RN(n2278), .QN(n1414)
         );
  DFFRXL \reg_file_reg[22][19]  ( .D(n1015), .CK(clk), .RN(n2275), .QN(n1413)
         );
  DFFRXL \reg_file_reg[22][18]  ( .D(n1016), .CK(clk), .RN(n2283), .QN(n1412)
         );
  DFFRXL \reg_file_reg[22][17]  ( .D(n1017), .CK(clk), .RN(n2275), .QN(n1411)
         );
  DFFRXL \reg_file_reg[22][16]  ( .D(n1018), .CK(clk), .RN(n2276), .QN(n1410)
         );
  DFFRXL \reg_file_reg[22][15]  ( .D(n1019), .CK(clk), .RN(n2276), .QN(n1409)
         );
  DFFRXL \reg_file_reg[22][14]  ( .D(n1020), .CK(clk), .RN(n2277), .QN(n1408)
         );
  DFFRXL \reg_file_reg[22][13]  ( .D(n1021), .CK(clk), .RN(n2277), .QN(n1407)
         );
  DFFRXL \reg_file_reg[22][12]  ( .D(n1022), .CK(clk), .RN(n2278), .QN(n1406)
         );
  DFFRXL \reg_file_reg[22][11]  ( .D(n1023), .CK(clk), .RN(n2279), .QN(n1405)
         );
  DFFRXL \reg_file_reg[22][10]  ( .D(n1024), .CK(clk), .RN(n2279), .QN(n1404)
         );
  DFFRXL \reg_file_reg[22][9]  ( .D(n1025), .CK(clk), .RN(n2280), .QN(n1403)
         );
  DFFRXL \reg_file_reg[22][8]  ( .D(n1026), .CK(clk), .RN(n2280), .QN(n1402)
         );
  DFFRXL \reg_file_reg[22][7]  ( .D(n1027), .CK(clk), .RN(n2281), .QN(n1401)
         );
  DFFRXL \reg_file_reg[22][6]  ( .D(n1028), .CK(clk), .RN(n2281), .QN(n1400)
         );
  DFFRXL \reg_file_reg[22][5]  ( .D(n1029), .CK(clk), .RN(n2283), .QN(n1399)
         );
  DFFRXL \reg_file_reg[22][4]  ( .D(n1030), .CK(clk), .RN(n2283), .QN(n1398)
         );
  DFFRXL \reg_file_reg[22][3]  ( .D(n1031), .CK(clk), .RN(n2282), .QN(n1397)
         );
  DFFRXL \reg_file_reg[22][2]  ( .D(n1032), .CK(clk), .RN(n2282), .QN(n1396)
         );
  DFFRXL \reg_file_reg[22][1]  ( .D(n1033), .CK(clk), .RN(n2282), .QN(n1395)
         );
  DFFRXL \reg_file_reg[22][0]  ( .D(n1034), .CK(clk), .RN(n2282), .QN(n1394)
         );
  DFFRXL \reg_file_reg[23][31]  ( .D(n1035), .CK(clk), .RN(n2284), .QN(n1393)
         );
  DFFRXL \reg_file_reg[23][30]  ( .D(n1036), .CK(clk), .RN(n2271), .QN(n1392)
         );
  DFFRXL \reg_file_reg[23][29]  ( .D(n1037), .CK(clk), .RN(n2271), .QN(n1391)
         );
  DFFRXL \reg_file_reg[23][28]  ( .D(n1038), .CK(clk), .RN(n2272), .QN(n1390)
         );
  DFFRXL \reg_file_reg[23][27]  ( .D(n1039), .CK(clk), .RN(n2272), .QN(n1389)
         );
  DFFRXL \reg_file_reg[23][26]  ( .D(n1040), .CK(clk), .RN(n2273), .QN(n1388)
         );
  DFFRXL \reg_file_reg[23][25]  ( .D(n1041), .CK(clk), .RN(n2273), .QN(n1387)
         );
  DFFRXL \reg_file_reg[23][24]  ( .D(n1042), .CK(clk), .RN(n2275), .QN(n1386)
         );
  DFFRXL \reg_file_reg[23][23]  ( .D(n1043), .CK(clk), .RN(n2274), .QN(n1385)
         );
  DFFRXL \reg_file_reg[23][22]  ( .D(n1044), .CK(clk), .RN(n2274), .QN(n1384)
         );
  DFFRXL \reg_file_reg[23][21]  ( .D(n1045), .CK(clk), .RN(n2279), .QN(n1383)
         );
  DFFRXL \reg_file_reg[23][20]  ( .D(n1046), .CK(clk), .RN(n2271), .QN(n1382)
         );
  DFFRXL \reg_file_reg[23][19]  ( .D(n1047), .CK(clk), .RN(n2275), .QN(n1381)
         );
  DFFRXL \reg_file_reg[23][18]  ( .D(n1048), .CK(clk), .RN(n2282), .QN(n1380)
         );
  DFFRXL \reg_file_reg[23][17]  ( .D(n1049), .CK(clk), .RN(n2275), .QN(n1379)
         );
  DFFRXL \reg_file_reg[23][16]  ( .D(n1050), .CK(clk), .RN(n2276), .QN(n1378)
         );
  DFFRXL \reg_file_reg[23][15]  ( .D(n1051), .CK(clk), .RN(n2276), .QN(n1377)
         );
  DFFRXL \reg_file_reg[23][14]  ( .D(n1052), .CK(clk), .RN(n2277), .QN(n1376)
         );
  DFFRXL \reg_file_reg[23][13]  ( .D(n1053), .CK(clk), .RN(n2277), .QN(n1375)
         );
  DFFRXL \reg_file_reg[23][12]  ( .D(n1054), .CK(clk), .RN(n2278), .QN(n1374)
         );
  DFFRXL \reg_file_reg[23][11]  ( .D(n1055), .CK(clk), .RN(n2279), .QN(n1373)
         );
  DFFRXL \reg_file_reg[23][10]  ( .D(n1056), .CK(clk), .RN(n2279), .QN(n1372)
         );
  DFFRXL \reg_file_reg[23][9]  ( .D(n1057), .CK(clk), .RN(n2280), .QN(n1371)
         );
  DFFRXL \reg_file_reg[23][8]  ( .D(n1058), .CK(clk), .RN(n2280), .QN(n1370)
         );
  DFFRXL \reg_file_reg[23][7]  ( .D(n1059), .CK(clk), .RN(n2281), .QN(n1369)
         );
  DFFRXL \reg_file_reg[23][6]  ( .D(n1060), .CK(clk), .RN(n2281), .QN(n1368)
         );
  DFFRXL \reg_file_reg[23][5]  ( .D(n1061), .CK(clk), .RN(n2282), .QN(n1367)
         );
  DFFRXL \reg_file_reg[23][4]  ( .D(n1062), .CK(clk), .RN(n2282), .QN(n1366)
         );
  DFFRXL \reg_file_reg[23][3]  ( .D(n1063), .CK(clk), .RN(n2282), .QN(n1365)
         );
  DFFRXL \reg_file_reg[23][2]  ( .D(n1064), .CK(clk), .RN(n2282), .QN(n1364)
         );
  DFFRXL \reg_file_reg[23][1]  ( .D(n1065), .CK(clk), .RN(n2282), .QN(n1363)
         );
  DFFRXL \reg_file_reg[23][0]  ( .D(n1066), .CK(clk), .RN(n2282), .QN(n1362)
         );
  DFFRXL \reg_file_reg[24][31]  ( .D(n1067), .CK(clk), .RN(n2283), .QN(n1361)
         );
  DFFRXL \reg_file_reg[24][30]  ( .D(n1068), .CK(clk), .RN(n2271), .QN(n1360)
         );
  DFFRXL \reg_file_reg[24][29]  ( .D(n1069), .CK(clk), .RN(n2271), .QN(n1359)
         );
  DFFRXL \reg_file_reg[24][28]  ( .D(n1070), .CK(clk), .RN(n2272), .QN(n1358)
         );
  DFFRXL \reg_file_reg[24][27]  ( .D(n1071), .CK(clk), .RN(n2272), .QN(n1357)
         );
  DFFRXL \reg_file_reg[24][26]  ( .D(n1072), .CK(clk), .RN(n2273), .QN(n1356)
         );
  DFFRXL \reg_file_reg[24][25]  ( .D(n1073), .CK(clk), .RN(n2273), .QN(n1355)
         );
  DFFRXL \reg_file_reg[24][24]  ( .D(n1074), .CK(clk), .RN(n2280), .QN(n298)
         );
  DFFRXL \reg_file_reg[24][23]  ( .D(n1075), .CK(clk), .RN(n2281), .QN(n297)
         );
  DFFRXL \reg_file_reg[24][22]  ( .D(n1076), .CK(clk), .RN(n2274), .QN(n296)
         );
  DFFRXL \reg_file_reg[24][21]  ( .D(n1077), .CK(clk), .RN(n2274), .QN(n295)
         );
  DFFRXL \reg_file_reg[24][20]  ( .D(n1078), .CK(clk), .RN(n2277), .QN(n294)
         );
  DFFRXL \reg_file_reg[24][19]  ( .D(n1079), .CK(clk), .RN(n2275), .QN(n293)
         );
  DFFRXL \reg_file_reg[24][18]  ( .D(n1080), .CK(clk), .RN(n2283), .QN(n292)
         );
  DFFRXL \reg_file_reg[24][17]  ( .D(n1081), .CK(clk), .RN(n2275), .QN(n291)
         );
  DFFRXL \reg_file_reg[24][16]  ( .D(n1082), .CK(clk), .RN(n2276), .QN(n290)
         );
  DFFRXL \reg_file_reg[24][15]  ( .D(n1083), .CK(clk), .RN(n2276), .QN(n289)
         );
  DFFRXL \reg_file_reg[24][14]  ( .D(n1084), .CK(clk), .RN(n2277), .QN(n288)
         );
  DFFRXL \reg_file_reg[24][13]  ( .D(n1085), .CK(clk), .RN(n2277), .QN(n287)
         );
  DFFRXL \reg_file_reg[24][12]  ( .D(n1086), .CK(clk), .RN(n2278), .QN(n286)
         );
  DFFRXL \reg_file_reg[24][11]  ( .D(n1087), .CK(clk), .RN(n2279), .QN(n285)
         );
  DFFRXL \reg_file_reg[24][10]  ( .D(n1088), .CK(clk), .RN(n2279), .QN(n284)
         );
  DFFRXL \reg_file_reg[24][9]  ( .D(n1089), .CK(clk), .RN(n2280), .QN(n283) );
  DFFRXL \reg_file_reg[24][8]  ( .D(n1090), .CK(clk), .RN(n2280), .QN(n282) );
  DFFRXL \reg_file_reg[24][7]  ( .D(n1091), .CK(clk), .RN(n2281), .QN(n281) );
  DFFRXL \reg_file_reg[24][6]  ( .D(n1092), .CK(clk), .RN(n2281), .QN(n280) );
  DFFRXL \reg_file_reg[24][5]  ( .D(n1093), .CK(clk), .RN(n2283), .QN(n279) );
  DFFRXL \reg_file_reg[24][4]  ( .D(n1094), .CK(clk), .RN(n2283), .QN(n278) );
  DFFRXL \reg_file_reg[24][3]  ( .D(n1095), .CK(clk), .RN(n2283), .QN(n277) );
  DFFRXL \reg_file_reg[24][2]  ( .D(n1096), .CK(clk), .RN(n2282), .QN(n276) );
  DFFRXL \reg_file_reg[24][1]  ( .D(n1097), .CK(clk), .RN(n2283), .QN(n275) );
  DFFRXL \reg_file_reg[24][0]  ( .D(n1098), .CK(clk), .RN(n2283), .QN(n274) );
  DFFRXL \reg_file_reg[25][31]  ( .D(n1099), .CK(clk), .RN(n2284), .QN(n273)
         );
  DFFRXL \reg_file_reg[25][30]  ( .D(n1100), .CK(clk), .RN(n2271), .QN(n272)
         );
  DFFRXL \reg_file_reg[25][29]  ( .D(n1101), .CK(clk), .RN(n2271), .QN(n271)
         );
  DFFRXL \reg_file_reg[25][28]  ( .D(n1102), .CK(clk), .RN(n2272), .QN(n270)
         );
  DFFRXL \reg_file_reg[25][27]  ( .D(n1103), .CK(clk), .RN(n2272), .QN(n269)
         );
  DFFRXL \reg_file_reg[25][26]  ( .D(n1104), .CK(clk), .RN(n2273), .QN(n268)
         );
  DFFRXL \reg_file_reg[25][25]  ( .D(n1105), .CK(clk), .RN(n2273), .QN(n267)
         );
  DFFRXL \reg_file_reg[25][24]  ( .D(n1106), .CK(clk), .RN(n2283), .QN(n266)
         );
  DFFRXL \reg_file_reg[25][23]  ( .D(n1107), .CK(clk), .RN(n2284), .QN(n265)
         );
  DFFRXL \reg_file_reg[25][22]  ( .D(n1108), .CK(clk), .RN(n2274), .QN(n264)
         );
  DFFRXL \reg_file_reg[25][21]  ( .D(n1109), .CK(clk), .RN(n2273), .QN(n263)
         );
  DFFRXL \reg_file_reg[25][20]  ( .D(n1110), .CK(clk), .RN(n2272), .QN(n262)
         );
  DFFRXL \reg_file_reg[25][19]  ( .D(n1111), .CK(clk), .RN(n2275), .QN(n261)
         );
  DFFRXL \reg_file_reg[25][18]  ( .D(n1112), .CK(clk), .RN(n2283), .QN(n260)
         );
  DFFRXL \reg_file_reg[25][17]  ( .D(n1113), .CK(clk), .RN(n2275), .QN(n259)
         );
  DFFRXL \reg_file_reg[25][16]  ( .D(n1114), .CK(clk), .RN(n2276), .QN(n258)
         );
  DFFRXL \reg_file_reg[25][15]  ( .D(n1115), .CK(clk), .RN(n2276), .QN(n257)
         );
  DFFRXL \reg_file_reg[25][14]  ( .D(n1116), .CK(clk), .RN(n2277), .QN(n256)
         );
  DFFRXL \reg_file_reg[25][13]  ( .D(n1117), .CK(clk), .RN(n2277), .QN(n255)
         );
  DFFRXL \reg_file_reg[25][12]  ( .D(n1118), .CK(clk), .RN(n2278), .QN(n254)
         );
  DFFRXL \reg_file_reg[25][11]  ( .D(n1119), .CK(clk), .RN(n2279), .QN(n253)
         );
  DFFRXL \reg_file_reg[25][10]  ( .D(n1120), .CK(clk), .RN(n2279), .QN(n252)
         );
  DFFRXL \reg_file_reg[25][9]  ( .D(n1121), .CK(clk), .RN(n2280), .QN(n251) );
  DFFRXL \reg_file_reg[25][8]  ( .D(n1122), .CK(clk), .RN(n2280), .QN(n250) );
  DFFRXL \reg_file_reg[25][7]  ( .D(n1123), .CK(clk), .RN(n2281), .QN(n249) );
  DFFRXL \reg_file_reg[25][6]  ( .D(n1124), .CK(clk), .RN(n2281), .QN(n248) );
  DFFRXL \reg_file_reg[25][5]  ( .D(n1125), .CK(clk), .RN(n2283), .QN(n247) );
  DFFRXL \reg_file_reg[25][4]  ( .D(n1126), .CK(clk), .RN(n2283), .QN(n246) );
  DFFRXL \reg_file_reg[25][3]  ( .D(n1127), .CK(clk), .RN(n2283), .QN(n245) );
  DFFRXL \reg_file_reg[25][2]  ( .D(n1128), .CK(clk), .RN(n2282), .QN(n244) );
  DFFRXL \reg_file_reg[25][1]  ( .D(n1129), .CK(clk), .RN(n2283), .QN(n243) );
  DFFRXL \reg_file_reg[25][0]  ( .D(n1130), .CK(clk), .RN(n2283), .QN(n242) );
  DFFRXL \reg_file_reg[26][31]  ( .D(n1131), .CK(clk), .RN(n2278), .QN(n241)
         );
  DFFRXL \reg_file_reg[26][30]  ( .D(n1132), .CK(clk), .RN(n2271), .QN(n240)
         );
  DFFRXL \reg_file_reg[26][29]  ( .D(n1133), .CK(clk), .RN(n2271), .QN(n239)
         );
  DFFRXL \reg_file_reg[26][28]  ( .D(n1134), .CK(clk), .RN(n2272), .QN(n238)
         );
  DFFRXL \reg_file_reg[26][27]  ( .D(n1135), .CK(clk), .RN(n2272), .QN(n237)
         );
  DFFRXL \reg_file_reg[26][26]  ( .D(n1136), .CK(clk), .RN(n2273), .QN(n236)
         );
  DFFRXL \reg_file_reg[26][25]  ( .D(n1137), .CK(clk), .RN(n2273), .QN(n235)
         );
  DFFRXL \reg_file_reg[26][24]  ( .D(n1138), .CK(clk), .RN(n2282), .QN(n234)
         );
  DFFRXL \reg_file_reg[26][23]  ( .D(n1139), .CK(clk), .RN(n2278), .QN(n233)
         );
  DFFRXL \reg_file_reg[26][22]  ( .D(n1140), .CK(clk), .RN(n2274), .QN(n232)
         );
  DFFRXL \reg_file_reg[26][21]  ( .D(n1141), .CK(clk), .RN(n2281), .QN(n231)
         );
  DFFRXL \reg_file_reg[26][20]  ( .D(n1142), .CK(clk), .RN(n2276), .QN(n230)
         );
  DFFRXL \reg_file_reg[26][19]  ( .D(n1143), .CK(clk), .RN(n2275), .QN(n229)
         );
  DFFRXL \reg_file_reg[26][18]  ( .D(n1144), .CK(clk), .RN(n2283), .QN(n228)
         );
  DFFRXL \reg_file_reg[26][17]  ( .D(n1145), .CK(clk), .RN(n2275), .QN(n227)
         );
  DFFRXL \reg_file_reg[26][16]  ( .D(n1146), .CK(clk), .RN(n2276), .QN(n226)
         );
  DFFRXL \reg_file_reg[26][15]  ( .D(n1147), .CK(clk), .RN(n2276), .QN(n225)
         );
  DFFRXL \reg_file_reg[26][14]  ( .D(n1148), .CK(clk), .RN(n2277), .QN(n224)
         );
  DFFRXL \reg_file_reg[26][13]  ( .D(n1149), .CK(clk), .RN(n2277), .QN(n223)
         );
  DFFRXL \reg_file_reg[26][12]  ( .D(n1150), .CK(clk), .RN(n2278), .QN(n222)
         );
  DFFRXL \reg_file_reg[26][11]  ( .D(n1151), .CK(clk), .RN(n2278), .QN(n221)
         );
  DFFRXL \reg_file_reg[26][10]  ( .D(n1152), .CK(clk), .RN(n2279), .QN(n220)
         );
  DFFRXL \reg_file_reg[26][9]  ( .D(n1153), .CK(clk), .RN(n2280), .QN(n219) );
  DFFRXL \reg_file_reg[26][8]  ( .D(n1154), .CK(clk), .RN(n2280), .QN(n218) );
  DFFRXL \reg_file_reg[26][7]  ( .D(n1155), .CK(clk), .RN(n2281), .QN(n217) );
  DFFRXL \reg_file_reg[26][6]  ( .D(n1156), .CK(clk), .RN(n2281), .QN(n216) );
  DFFRXL \reg_file_reg[26][5]  ( .D(n1157), .CK(clk), .RN(n2283), .QN(n215) );
  DFFRXL \reg_file_reg[26][4]  ( .D(n1158), .CK(clk), .RN(n2283), .QN(n214) );
  DFFRXL \reg_file_reg[26][3]  ( .D(n1159), .CK(clk), .RN(n2283), .QN(n213) );
  DFFRXL \reg_file_reg[26][2]  ( .D(n1160), .CK(clk), .RN(n2282), .QN(n212) );
  DFFRXL \reg_file_reg[26][1]  ( .D(n1161), .CK(clk), .RN(n2283), .QN(n211) );
  DFFRXL \reg_file_reg[26][0]  ( .D(n1162), .CK(clk), .RN(n2283), .QN(n210) );
  DFFRXL \reg_file_reg[27][31]  ( .D(n1163), .CK(clk), .RN(n2282), .QN(n209)
         );
  DFFRXL \reg_file_reg[27][30]  ( .D(n1164), .CK(clk), .RN(n2271), .QN(n208)
         );
  DFFRXL \reg_file_reg[27][29]  ( .D(n1165), .CK(clk), .RN(n2271), .QN(n207)
         );
  DFFRXL \reg_file_reg[27][28]  ( .D(n1166), .CK(clk), .RN(n2272), .QN(n206)
         );
  DFFRXL \reg_file_reg[27][27]  ( .D(n1167), .CK(clk), .RN(n2272), .QN(n205)
         );
  DFFRXL \reg_file_reg[27][26]  ( .D(n1168), .CK(clk), .RN(n2273), .QN(n204)
         );
  DFFRXL \reg_file_reg[27][25]  ( .D(n1169), .CK(clk), .RN(n2273), .QN(n203)
         );
  DFFRXL \reg_file_reg[27][24]  ( .D(n1170), .CK(clk), .RN(n2279), .QN(n202)
         );
  DFFRXL \reg_file_reg[27][23]  ( .D(n1171), .CK(clk), .RN(n2271), .QN(n201)
         );
  DFFRXL \reg_file_reg[27][22]  ( .D(n1172), .CK(clk), .RN(n2274), .QN(n200)
         );
  DFFRXL \reg_file_reg[27][21]  ( .D(n1173), .CK(clk), .RN(n2275), .QN(n199)
         );
  DFFRXL \reg_file_reg[27][20]  ( .D(n1174), .CK(clk), .RN(n2280), .QN(n198)
         );
  DFFRXL \reg_file_reg[27][19]  ( .D(n1175), .CK(clk), .RN(n2275), .QN(n197)
         );
  DFFRXL \reg_file_reg[27][18]  ( .D(n1176), .CK(clk), .RN(n2283), .QN(n196)
         );
  DFFRXL \reg_file_reg[27][17]  ( .D(n1177), .CK(clk), .RN(n2275), .QN(n195)
         );
  DFFRXL \reg_file_reg[27][16]  ( .D(n1178), .CK(clk), .RN(n2276), .QN(n194)
         );
  DFFRXL \reg_file_reg[27][15]  ( .D(n1179), .CK(clk), .RN(n2276), .QN(n193)
         );
  DFFRXL \reg_file_reg[27][14]  ( .D(n1180), .CK(clk), .RN(n2277), .QN(n192)
         );
  DFFRXL \reg_file_reg[27][13]  ( .D(n1181), .CK(clk), .RN(n2277), .QN(n191)
         );
  DFFRXL \reg_file_reg[27][12]  ( .D(n1182), .CK(clk), .RN(n2278), .QN(n190)
         );
  DFFRXL \reg_file_reg[27][11]  ( .D(n1183), .CK(clk), .RN(n2278), .QN(n189)
         );
  DFFRXL \reg_file_reg[27][10]  ( .D(n1184), .CK(clk), .RN(n2279), .QN(n188)
         );
  DFFRXL \reg_file_reg[27][9]  ( .D(n1185), .CK(clk), .RN(n2280), .QN(n187) );
  DFFRXL \reg_file_reg[27][8]  ( .D(n1186), .CK(clk), .RN(n2280), .QN(n186) );
  DFFRXL \reg_file_reg[27][7]  ( .D(n1187), .CK(clk), .RN(n2281), .QN(n185) );
  DFFRXL \reg_file_reg[27][6]  ( .D(n1188), .CK(clk), .RN(n2281), .QN(n184) );
  DFFRXL \reg_file_reg[27][5]  ( .D(n1189), .CK(clk), .RN(n2283), .QN(n183) );
  DFFRXL \reg_file_reg[27][4]  ( .D(n1190), .CK(clk), .RN(n2283), .QN(n182) );
  DFFRXL \reg_file_reg[27][3]  ( .D(n1191), .CK(clk), .RN(n2283), .QN(n181) );
  DFFRXL \reg_file_reg[27][2]  ( .D(n1192), .CK(clk), .RN(n2282), .QN(n180) );
  DFFRXL \reg_file_reg[27][1]  ( .D(n1193), .CK(clk), .RN(n2283), .QN(n179) );
  DFFRXL \reg_file_reg[27][0]  ( .D(n1194), .CK(clk), .RN(n2283), .QN(n178) );
  DFFRXL \reg_file_reg[28][31]  ( .D(n1195), .CK(clk), .RN(n2285), .QN(n177)
         );
  DFFRXL \reg_file_reg[28][30]  ( .D(n1196), .CK(clk), .RN(n2271), .QN(n176)
         );
  DFFRXL \reg_file_reg[28][29]  ( .D(n1197), .CK(clk), .RN(n2271), .QN(n175)
         );
  DFFRXL \reg_file_reg[28][28]  ( .D(n1198), .CK(clk), .RN(n2272), .QN(n174)
         );
  DFFRXL \reg_file_reg[28][27]  ( .D(n1199), .CK(clk), .RN(n2272), .QN(n173)
         );
  DFFRXL \reg_file_reg[28][26]  ( .D(n1200), .CK(clk), .RN(n2273), .QN(n172)
         );
  DFFRXL \reg_file_reg[28][25]  ( .D(n1201), .CK(clk), .RN(n2273), .QN(n171)
         );
  DFFRXL \reg_file_reg[28][24]  ( .D(n1202), .CK(clk), .RN(n2274), .QN(n170)
         );
  DFFRXL \reg_file_reg[28][23]  ( .D(n1203), .CK(clk), .RN(n2277), .QN(n169)
         );
  DFFRXL \reg_file_reg[28][22]  ( .D(n1204), .CK(clk), .RN(n2274), .QN(n168)
         );
  DFFRXL \reg_file_reg[28][21]  ( .D(n1205), .CK(clk), .RN(n2283), .QN(n167)
         );
  DFFRXL \reg_file_reg[28][20]  ( .D(n1206), .CK(clk), .RN(n2284), .QN(n166)
         );
  DFFRXL \reg_file_reg[28][19]  ( .D(n1207), .CK(clk), .RN(n2275), .QN(n165)
         );
  DFFRXL \reg_file_reg[28][18]  ( .D(n1208), .CK(clk), .RN(n2283), .QN(n164)
         );
  DFFRXL \reg_file_reg[28][17]  ( .D(n1209), .CK(clk), .RN(n2275), .QN(n163)
         );
  DFFRXL \reg_file_reg[28][16]  ( .D(n1210), .CK(clk), .RN(n2276), .QN(n162)
         );
  DFFRXL \reg_file_reg[28][15]  ( .D(n1211), .CK(clk), .RN(n2276), .QN(n161)
         );
  DFFRXL \reg_file_reg[28][14]  ( .D(n1212), .CK(clk), .RN(n2277), .QN(n160)
         );
  DFFRXL \reg_file_reg[28][13]  ( .D(n1213), .CK(clk), .RN(n2277), .QN(n159)
         );
  DFFRXL \reg_file_reg[28][12]  ( .D(n1214), .CK(clk), .RN(n2278), .QN(n158)
         );
  DFFRXL \reg_file_reg[28][11]  ( .D(n1215), .CK(clk), .RN(n2278), .QN(n157)
         );
  DFFRXL \reg_file_reg[28][10]  ( .D(n1216), .CK(clk), .RN(n2279), .QN(n156)
         );
  DFFRXL \reg_file_reg[28][9]  ( .D(n1217), .CK(clk), .RN(n2280), .QN(n155) );
  DFFRXL \reg_file_reg[28][8]  ( .D(n1218), .CK(clk), .RN(n2280), .QN(n154) );
  DFFRXL \reg_file_reg[28][7]  ( .D(n1219), .CK(clk), .RN(n2281), .QN(n153) );
  DFFRXL \reg_file_reg[28][6]  ( .D(n1220), .CK(clk), .RN(n2281), .QN(n152) );
  DFFRXL \reg_file_reg[28][5]  ( .D(n1221), .CK(clk), .RN(n2283), .QN(n151) );
  DFFRXL \reg_file_reg[28][4]  ( .D(n1222), .CK(clk), .RN(n2283), .QN(n150) );
  DFFRXL \reg_file_reg[28][3]  ( .D(n1223), .CK(clk), .RN(n2283), .QN(n149) );
  DFFRXL \reg_file_reg[28][2]  ( .D(n1224), .CK(clk), .RN(n2282), .QN(n148) );
  DFFRXL \reg_file_reg[28][1]  ( .D(n1225), .CK(clk), .RN(n2283), .QN(n147) );
  DFFRXL \reg_file_reg[28][0]  ( .D(n1226), .CK(clk), .RN(n2283), .QN(n146) );
  DFFRXL \reg_file_reg[29][31]  ( .D(n1227), .CK(clk), .RN(n2285), .QN(n145)
         );
  DFFRXL \reg_file_reg[29][30]  ( .D(n1228), .CK(clk), .RN(n2271), .QN(n144)
         );
  DFFRXL \reg_file_reg[29][29]  ( .D(n1229), .CK(clk), .RN(n2271), .QN(n143)
         );
  DFFRXL \reg_file_reg[29][28]  ( .D(n1230), .CK(clk), .RN(n2272), .QN(n142)
         );
  DFFRXL \reg_file_reg[29][27]  ( .D(n1231), .CK(clk), .RN(n2272), .QN(n141)
         );
  DFFRXL \reg_file_reg[29][26]  ( .D(n1232), .CK(clk), .RN(n2273), .QN(n140)
         );
  DFFRXL \reg_file_reg[29][25]  ( .D(n1233), .CK(clk), .RN(n2273), .QN(n139)
         );
  DFFRXL \reg_file_reg[29][24]  ( .D(n1234), .CK(clk), .RN(n2273), .QN(n138)
         );
  DFFRXL \reg_file_reg[29][23]  ( .D(n1235), .CK(clk), .RN(n2272), .QN(n137)
         );
  DFFRXL \reg_file_reg[29][22]  ( .D(n1236), .CK(clk), .RN(n2274), .QN(n136)
         );
  DFFRXL \reg_file_reg[29][21]  ( .D(n1237), .CK(clk), .RN(n2282), .QN(n135)
         );
  DFFRXL \reg_file_reg[29][20]  ( .D(n1238), .CK(clk), .RN(n2278), .QN(n134)
         );
  DFFRXL \reg_file_reg[29][19]  ( .D(n1239), .CK(clk), .RN(n2275), .QN(n133)
         );
  DFFRXL \reg_file_reg[29][18]  ( .D(n1240), .CK(clk), .RN(n2283), .QN(n132)
         );
  DFFRXL \reg_file_reg[29][17]  ( .D(n1241), .CK(clk), .RN(n2275), .QN(n131)
         );
  DFFRXL \reg_file_reg[29][16]  ( .D(n1242), .CK(clk), .RN(n2276), .QN(n130)
         );
  DFFRXL \reg_file_reg[29][15]  ( .D(n1243), .CK(clk), .RN(n2276), .QN(n129)
         );
  DFFRXL \reg_file_reg[29][14]  ( .D(n1244), .CK(clk), .RN(n2277), .QN(n128)
         );
  DFFRXL \reg_file_reg[29][13]  ( .D(n1245), .CK(clk), .RN(n2277), .QN(n127)
         );
  DFFRXL \reg_file_reg[29][12]  ( .D(n1246), .CK(clk), .RN(n2278), .QN(n126)
         );
  DFFRXL \reg_file_reg[29][11]  ( .D(n1247), .CK(clk), .RN(n2278), .QN(n125)
         );
  DFFRXL \reg_file_reg[29][10]  ( .D(n1248), .CK(clk), .RN(n2279), .QN(n124)
         );
  DFFRXL \reg_file_reg[29][9]  ( .D(n1249), .CK(clk), .RN(n2280), .QN(n123) );
  DFFRXL \reg_file_reg[29][8]  ( .D(n1250), .CK(clk), .RN(n2280), .QN(n122) );
  DFFRXL \reg_file_reg[29][7]  ( .D(n1251), .CK(clk), .RN(n2281), .QN(n121) );
  DFFRXL \reg_file_reg[29][6]  ( .D(n1252), .CK(clk), .RN(n2281), .QN(n120) );
  DFFRXL \reg_file_reg[29][5]  ( .D(n1253), .CK(clk), .RN(n2283), .QN(n119) );
  DFFRXL \reg_file_reg[29][4]  ( .D(n1254), .CK(clk), .RN(n2283), .QN(n118) );
  DFFRXL \reg_file_reg[29][3]  ( .D(n1255), .CK(clk), .RN(n2283), .QN(n117) );
  DFFRXL \reg_file_reg[29][2]  ( .D(n1256), .CK(clk), .RN(n2282), .QN(n116) );
  DFFRXL \reg_file_reg[29][1]  ( .D(n1257), .CK(clk), .RN(n2283), .QN(n115) );
  DFFRXL \reg_file_reg[29][0]  ( .D(n1258), .CK(clk), .RN(n2283), .QN(n114) );
  DFFRXL \reg_file_reg[30][31]  ( .D(n1259), .CK(clk), .RN(n2285), .QN(n113)
         );
  DFFRXL \reg_file_reg[30][30]  ( .D(n1260), .CK(clk), .RN(n2271), .QN(n112)
         );
  DFFRXL \reg_file_reg[30][29]  ( .D(n1261), .CK(clk), .RN(n2271), .QN(n111)
         );
  DFFRXL \reg_file_reg[30][28]  ( .D(n1262), .CK(clk), .RN(n2272), .QN(n110)
         );
  DFFRXL \reg_file_reg[30][27]  ( .D(n1263), .CK(clk), .RN(n2272), .QN(n109)
         );
  DFFRXL \reg_file_reg[30][26]  ( .D(n1264), .CK(clk), .RN(n2273), .QN(n108)
         );
  DFFRXL \reg_file_reg[30][25]  ( .D(n1265), .CK(clk), .RN(n2273), .QN(n107)
         );
  DFFRXL \reg_file_reg[30][24]  ( .D(n1266), .CK(clk), .RN(n2276), .QN(n106)
         );
  DFFRXL \reg_file_reg[30][23]  ( .D(n1267), .CK(clk), .RN(n2280), .QN(n105)
         );
  DFFRXL \reg_file_reg[30][22]  ( .D(n1268), .CK(clk), .RN(n2274), .QN(n104)
         );
  DFFRXL \reg_file_reg[30][21]  ( .D(n1269), .CK(clk), .RN(n2274), .QN(n103)
         );
  DFFRXL \reg_file_reg[30][20]  ( .D(n1270), .CK(clk), .RN(n2279), .QN(n102)
         );
  DFFRXL \reg_file_reg[30][19]  ( .D(n1271), .CK(clk), .RN(n2275), .QN(n101)
         );
  DFFRXL \reg_file_reg[30][18]  ( .D(n1272), .CK(clk), .RN(n2283), .QN(n100)
         );
  DFFRXL \reg_file_reg[30][17]  ( .D(n1273), .CK(clk), .RN(n2275), .QN(n99) );
  DFFRXL \reg_file_reg[30][16]  ( .D(n1274), .CK(clk), .RN(n2276), .QN(n98) );
  DFFRXL \reg_file_reg[30][15]  ( .D(n1275), .CK(clk), .RN(n2276), .QN(n97) );
  DFFRXL \reg_file_reg[30][14]  ( .D(n1276), .CK(clk), .RN(n2277), .QN(n96) );
  DFFRXL \reg_file_reg[30][13]  ( .D(n1277), .CK(clk), .RN(n2277), .QN(n95) );
  DFFRXL \reg_file_reg[30][12]  ( .D(n1278), .CK(clk), .RN(n2278), .QN(n94) );
  DFFRXL \reg_file_reg[30][11]  ( .D(n1279), .CK(clk), .RN(n2278), .QN(n93) );
  DFFRXL \reg_file_reg[30][10]  ( .D(n1280), .CK(clk), .RN(n2279), .QN(n92) );
  DFFRXL \reg_file_reg[30][9]  ( .D(n1281), .CK(clk), .RN(n2280), .QN(n91) );
  DFFRXL \reg_file_reg[30][8]  ( .D(n1282), .CK(clk), .RN(n2280), .QN(n90) );
  DFFRXL \reg_file_reg[30][7]  ( .D(n1283), .CK(clk), .RN(n2281), .QN(n89) );
  DFFRXL \reg_file_reg[30][6]  ( .D(n1284), .CK(clk), .RN(n2281), .QN(n88) );
  DFFRXL \reg_file_reg[30][5]  ( .D(n1285), .CK(clk), .RN(n2283), .QN(n87) );
  DFFRXL \reg_file_reg[30][4]  ( .D(n1286), .CK(clk), .RN(n2283), .QN(n86) );
  DFFRXL \reg_file_reg[30][3]  ( .D(n1287), .CK(clk), .RN(n2283), .QN(n85) );
  DFFRXL \reg_file_reg[30][2]  ( .D(n1288), .CK(clk), .RN(n2282), .QN(n84) );
  DFFRXL \reg_file_reg[30][1]  ( .D(n1289), .CK(clk), .RN(n2283), .QN(n83) );
  DFFRXL \reg_file_reg[30][0]  ( .D(n1290), .CK(clk), .RN(n2283), .QN(n82) );
  DFFRXL \reg_file_reg[31][31]  ( .D(n1291), .CK(clk), .RN(n2285), .QN(n81) );
  DFFRXL \reg_file_reg[31][30]  ( .D(n1292), .CK(clk), .RN(n2271), .QN(n80) );
  DFFRXL \reg_file_reg[31][29]  ( .D(n1293), .CK(clk), .RN(n2271), .QN(n79) );
  DFFRXL \reg_file_reg[31][28]  ( .D(n1294), .CK(clk), .RN(n2272), .QN(n78) );
  DFFRXL \reg_file_reg[31][27]  ( .D(n1295), .CK(clk), .RN(n2272), .QN(n77) );
  DFFRXL \reg_file_reg[31][26]  ( .D(n1296), .CK(clk), .RN(n2273), .QN(n76) );
  DFFRXL \reg_file_reg[31][25]  ( .D(n1297), .CK(clk), .RN(n2273), .QN(n75) );
  DFFRXL \reg_file_reg[31][24]  ( .D(n1298), .CK(clk), .RN(n2275), .QN(n74) );
  DFFRXL \reg_file_reg[31][23]  ( .D(n1299), .CK(clk), .RN(n2280), .QN(n73) );
  DFFRXL \reg_file_reg[31][22]  ( .D(n1300), .CK(clk), .RN(n2274), .QN(n72) );
  DFFRXL \reg_file_reg[31][21]  ( .D(n1301), .CK(clk), .RN(n2274), .QN(n71) );
  DFFRXL \reg_file_reg[31][20]  ( .D(n1302), .CK(clk), .RN(n2271), .QN(n69) );
  DFFRXL \reg_file_reg[31][19]  ( .D(n1303), .CK(clk), .RN(n2275), .QN(n68) );
  DFFRXL \reg_file_reg[31][18]  ( .D(n1304), .CK(clk), .RN(n2283), .QN(n67) );
  DFFRXL \reg_file_reg[31][17]  ( .D(n1305), .CK(clk), .RN(n2275), .QN(n66) );
  DFFRXL \reg_file_reg[31][16]  ( .D(n1306), .CK(clk), .RN(n2276), .QN(n65) );
  DFFRXL \reg_file_reg[31][15]  ( .D(n1307), .CK(clk), .RN(n2276), .QN(n64) );
  DFFRXL \reg_file_reg[31][14]  ( .D(n1308), .CK(clk), .RN(n2277), .QN(n63) );
  DFFRXL \reg_file_reg[31][13]  ( .D(n1309), .CK(clk), .RN(n2277), .QN(n62) );
  DFFRXL \reg_file_reg[31][12]  ( .D(n1310), .CK(clk), .RN(n2278), .QN(n61) );
  DFFRXL \reg_file_reg[31][11]  ( .D(n1311), .CK(clk), .RN(n2278), .QN(n60) );
  DFFRXL \reg_file_reg[31][10]  ( .D(n1312), .CK(clk), .RN(n2279), .QN(n59) );
  DFFRXL \reg_file_reg[31][9]  ( .D(n1313), .CK(clk), .RN(n2280), .QN(n58) );
  DFFRXL \reg_file_reg[31][8]  ( .D(n1314), .CK(clk), .RN(n2280), .QN(n57) );
  DFFRXL \reg_file_reg[31][7]  ( .D(n1315), .CK(clk), .RN(n2281), .QN(n56) );
  DFFRXL \reg_file_reg[31][6]  ( .D(n1316), .CK(clk), .RN(n2281), .QN(n55) );
  DFFRXL \reg_file_reg[31][5]  ( .D(n1317), .CK(clk), .RN(n2283), .QN(n54) );
  DFFRXL \reg_file_reg[31][4]  ( .D(n1318), .CK(clk), .RN(n2283), .QN(n53) );
  DFFRXL \reg_file_reg[31][3]  ( .D(n1319), .CK(clk), .RN(n2283), .QN(n52) );
  DFFRXL \reg_file_reg[31][2]  ( .D(n1320), .CK(clk), .RN(n2282), .QN(n51) );
  DFFRXL \reg_file_reg[31][1]  ( .D(n1321), .CK(clk), .RN(n2283), .QN(n50) );
  DFFRXL \reg_file_reg[31][0]  ( .D(n1322), .CK(clk), .RN(n2283), .QN(n49) );
  DFFRX1 \IR_addr_reg[31]  ( .D(n1323), .CK(clk), .RN(n2285), .Q(
        ICACHE_addr[29]), .QN(n3220) );
  DFFRX1 \IR_addr_reg[10]  ( .D(n1344), .CK(clk), .RN(n2279), .Q(
        ICACHE_addr[8]), .QN(n3241) );
  DFFRX1 \IR_addr_reg[11]  ( .D(n1343), .CK(clk), .RN(n2279), .Q(
        ICACHE_addr[9]), .QN(n3240) );
  DFFRX1 \IR_addr_reg[12]  ( .D(n1342), .CK(clk), .RN(n2277), .Q(
        ICACHE_addr[10]), .QN(n3239) );
  DFFRX1 \IR_addr_reg[16]  ( .D(n1338), .CK(clk), .RN(n2275), .Q(
        ICACHE_addr[14]), .QN(n3235) );
  DFFRX1 \IR_addr_reg[17]  ( .D(n1337), .CK(clk), .RN(n2275), .Q(
        ICACHE_addr[15]), .QN(n3234) );
  DFFRX1 \IR_addr_reg[18]  ( .D(n1336), .CK(clk), .RN(n2285), .Q(
        ICACHE_addr[16]), .QN(n3233) );
  DFFRX1 \IR_addr_reg[22]  ( .D(n1332), .CK(clk), .RN(n2274), .Q(
        ICACHE_addr[20]), .QN(n3229) );
  DFFRX1 \IR_addr_reg[23]  ( .D(n1331), .CK(clk), .RN(rst_n), .Q(
        ICACHE_addr[21]), .QN(n3228) );
  DFFRX1 \IR_addr_reg[24]  ( .D(n1330), .CK(clk), .RN(n2273), .Q(
        ICACHE_addr[22]), .QN(n3227) );
  DFFRX1 \IR_addr_reg[28]  ( .D(n1326), .CK(clk), .RN(n2271), .Q(
        ICACHE_addr[26]), .QN(n3223) );
  DFFRX1 \IR_addr_reg[29]  ( .D(n1325), .CK(clk), .RN(n2271), .Q(
        ICACHE_addr[27]), .QN(n3222) );
  DFFRX1 \IR_addr_reg[30]  ( .D(n1324), .CK(clk), .RN(n2286), .Q(
        ICACHE_addr[28]), .QN(n3221) );
  DFFRX1 \IR_addr_reg[7]  ( .D(n1347), .CK(clk), .RN(n2281), .Q(ICACHE_addr[5]), .QN(n3244) );
  DFFRX1 \IR_addr_reg[8]  ( .D(n1346), .CK(clk), .RN(n2280), .Q(ICACHE_addr[6]), .QN(n3243) );
  DFFRX1 \IR_addr_reg[9]  ( .D(n1345), .CK(clk), .RN(n2280), .Q(ICACHE_addr[7]), .QN(n3242) );
  DFFRX1 \IR_addr_reg[13]  ( .D(n1341), .CK(clk), .RN(n2277), .Q(
        ICACHE_addr[11]), .QN(n3238) );
  DFFRX1 \IR_addr_reg[14]  ( .D(n1340), .CK(clk), .RN(n2276), .Q(
        ICACHE_addr[12]), .QN(n3237) );
  DFFRX1 \IR_addr_reg[15]  ( .D(n1339), .CK(clk), .RN(n2276), .Q(
        ICACHE_addr[13]), .QN(n3236) );
  DFFRX1 \IR_addr_reg[19]  ( .D(n1335), .CK(clk), .RN(n2281), .Q(
        ICACHE_addr[17]), .QN(n3232) );
  DFFRX1 \IR_addr_reg[20]  ( .D(n1334), .CK(clk), .RN(rst_n), .Q(
        ICACHE_addr[18]), .QN(n3231) );
  DFFRX1 \IR_addr_reg[21]  ( .D(n1333), .CK(clk), .RN(n2274), .Q(
        ICACHE_addr[19]), .QN(n3230) );
  DFFRX1 \IR_addr_reg[25]  ( .D(n1329), .CK(clk), .RN(n2273), .Q(
        ICACHE_addr[23]), .QN(n3226) );
  DFFRX1 \IR_addr_reg[26]  ( .D(n1328), .CK(clk), .RN(n2272), .Q(
        ICACHE_addr[24]), .QN(n3225) );
  DFFRX1 \IR_addr_reg[27]  ( .D(n1327), .CK(clk), .RN(n2272), .Q(
        ICACHE_addr[25]), .QN(n3224) );
  DFFRX2 \IR_addr_reg[2]  ( .D(n1352), .CK(clk), .RN(n2285), .Q(ICACHE_addr[0]), .QN(n3249) );
  DFFRXL \IR_addr_reg[4]  ( .D(n1350), .CK(clk), .RN(n2285), .Q(ICACHE_addr[2]), .QN(n3247) );
  DFFRXL \IR_addr_reg[5]  ( .D(n1349), .CK(clk), .RN(n2285), .Q(ICACHE_addr[3]), .QN(n3246) );
  DFFRX1 \IR_addr_reg[6]  ( .D(n1348), .CK(clk), .RN(n2285), .Q(ICACHE_addr[4]), .QN(n3245) );
  DFFRX4 \IR_addr_reg[3]  ( .D(n1351), .CK(clk), .RN(n2285), .Q(ICACHE_addr[1]), .QN(n3248) );
  OAI211X1 U40 ( .A0(n3245), .A1(n2139), .B0(n3047), .C0(n3048), .Y(n1348) );
  OR2X1 U41 ( .A(n3116), .B(ICACHE_stall), .Y(n43) );
  NAND3X1 U42 ( .A(Jump[0]), .B(n2139), .C(Jump[1]), .Y(n44) );
  AOI21X1 U43 ( .A0(M[0]), .A1(N1140), .B0(Jump[1]), .Y(n45) );
  XOR2X1 U44 ( .A(Foward_A[0]), .B(Foward_A[1]), .Y(n46) );
  XOR2X1 U45 ( .A(Foward_B[0]), .B(Foward_B[1]), .Y(n47) );
  NAND3X1 U46 ( .A(n3099), .B(n2139), .C(Jump[1]), .Y(n48) );
  INVXL U47 ( .A(n3249), .Y(n2130) );
  OAI21X2 U48 ( .A0(n3165), .A1(n2136), .B0(n3166), .Y(after_A_mux[17]) );
  OAI21X2 U49 ( .A0(n3123), .A1(n2136), .B0(n3124), .Y(after_A_mux[7]) );
  OAI21X2 U50 ( .A0(n3129), .A1(n2136), .B0(n3130), .Y(after_A_mux[4]) );
  OAI21X2 U51 ( .A0(n3135), .A1(n2136), .B0(n3136), .Y(after_A_mux[30]) );
  OAI21X2 U52 ( .A0(n3147), .A1(n2136), .B0(n3148), .Y(after_A_mux[25]) );
  OAI21X2 U53 ( .A0(n3181), .A1(n2136), .B0(n3182), .Y(after_A_mux[0]) );
  INVX8 U54 ( .A(n2135), .Y(n2136) );
  OAI21X2 U55 ( .A0(n3133), .A1(n2136), .B0(n3134), .Y(after_A_mux[31]) );
  OAI21X2 U56 ( .A0(n3167), .A1(n2136), .B0(n3168), .Y(after_A_mux[16]) );
  OAI21X2 U57 ( .A0(n3125), .A1(n2136), .B0(n3126), .Y(after_A_mux[6]) );
  OAI21X2 U58 ( .A0(n3149), .A1(n2136), .B0(n3150), .Y(after_A_mux[24]) );
  OAI21X2 U59 ( .A0(n3171), .A1(n2136), .B0(n3172), .Y(after_A_mux[14]) );
  OAI21X2 U60 ( .A0(n3153), .A1(n2136), .B0(n3154), .Y(after_A_mux[22]) );
  OAI21X2 U61 ( .A0(n3117), .A1(n2136), .B0(n3119), .Y(after_A_mux[9]) );
  OAI21X2 U62 ( .A0(n3157), .A1(n2136), .B0(n3158), .Y(after_A_mux[20]) );
  OAI21X2 U63 ( .A0(n3175), .A1(n2136), .B0(n3176), .Y(after_A_mux[12]) );
  OAI21X2 U64 ( .A0(n3137), .A1(n2136), .B0(n3138), .Y(after_A_mux[2]) );
  OAI21X2 U65 ( .A0(n3141), .A1(n2136), .B0(n3142), .Y(after_A_mux[28]) );
  OAI21X2 U66 ( .A0(n3163), .A1(n2136), .B0(n3164), .Y(after_A_mux[18]) );
  OAI21X2 U67 ( .A0(n3159), .A1(n2136), .B0(n3160), .Y(after_A_mux[1]) );
  OAI21X2 U68 ( .A0(n3177), .A1(n2136), .B0(n3178), .Y(after_A_mux[11]) );
  OAI21X2 U69 ( .A0(n3145), .A1(n2136), .B0(n3146), .Y(after_A_mux[26]) );
  OAI21X2 U70 ( .A0(n3169), .A1(n2136), .B0(n3170), .Y(after_A_mux[15]) );
  OAI21X2 U71 ( .A0(n3139), .A1(n2136), .B0(n3140), .Y(after_A_mux[29]) );
  OAI21X2 U72 ( .A0(n3127), .A1(n2136), .B0(n3128), .Y(after_A_mux[5]) );
  OAI21X2 U73 ( .A0(n3151), .A1(n2136), .B0(n3152), .Y(after_A_mux[23]) );
  OAI21X2 U74 ( .A0(n3161), .A1(n2136), .B0(n3162), .Y(after_A_mux[19]) );
  OAI21X2 U75 ( .A0(n3155), .A1(n2136), .B0(n3156), .Y(after_A_mux[21]) );
  OAI21X2 U76 ( .A0(n3173), .A1(n2136), .B0(n3174), .Y(after_A_mux[13]) );
  OAI21X2 U77 ( .A0(n3179), .A1(n2136), .B0(n3180), .Y(after_A_mux[10]) );
  OAI21X2 U78 ( .A0(n3131), .A1(n2136), .B0(n3132), .Y(after_A_mux[3]) );
  OAI21X2 U79 ( .A0(n3121), .A1(n2136), .B0(n3122), .Y(after_A_mux[8]) );
  OAI21X2 U80 ( .A0(n3143), .A1(n2136), .B0(n3144), .Y(after_A_mux[27]) );
  INVX6 U81 ( .A(n48), .Y(n2131) );
  CLKAND2X6 U82 ( .A(n2139), .B(n3100), .Y(n3035) );
  INVX6 U83 ( .A(n44), .Y(n2132) );
  CLKAND2X6 U84 ( .A(n2139), .B(n2966), .Y(n3102) );
  CLKAND2X6 U85 ( .A(n2139), .B(n2967), .Y(n3104) );
  CLKAND2X6 U86 ( .A(n2139), .B(n2969), .Y(n3105) );
  CLKAND2X6 U87 ( .A(n2139), .B(n2970), .Y(n3106) );
  CLKAND2X6 U88 ( .A(n2139), .B(n2971), .Y(n3108) );
  CLKAND2X6 U89 ( .A(n2139), .B(n2972), .Y(n3111) );
  CLKAND2X6 U90 ( .A(n2139), .B(n2973), .Y(n3112) );
  CLKAND2X6 U91 ( .A(n2139), .B(n2974), .Y(n3113) );
  CLKAND2X6 U92 ( .A(n2139), .B(n2975), .Y(n3114) );
  CLKAND2X6 U93 ( .A(n2139), .B(n2976), .Y(n3115) );
  CLKAND2X6 U94 ( .A(n2139), .B(n2977), .Y(n2991) );
  CLKAND2X6 U95 ( .A(n2139), .B(n2978), .Y(n2992) );
  CLKAND2X6 U96 ( .A(n2139), .B(n2980), .Y(n2995) );
  CLKAND2X6 U97 ( .A(n2139), .B(n2981), .Y(n2997) );
  CLKAND2X6 U98 ( .A(n2139), .B(n2982), .Y(n2999) );
  CLKAND2X6 U99 ( .A(n2139), .B(n2983), .Y(n3001) );
  CLKAND2X6 U100 ( .A(n2139), .B(n2984), .Y(n3003) );
  CLKAND2X6 U101 ( .A(n2139), .B(n2985), .Y(n3006) );
  CLKAND2X6 U102 ( .A(n2139), .B(n2986), .Y(n3008) );
  CLKAND2X6 U103 ( .A(n2139), .B(n2987), .Y(n3010) );
  CLKAND2X6 U104 ( .A(n2139), .B(n2988), .Y(n3011) );
  CLKAND2X6 U105 ( .A(n2139), .B(n2989), .Y(n3012) );
  CLKAND2X6 U106 ( .A(n2139), .B(n2928), .Y(n3013) );
  CLKAND2X6 U107 ( .A(n2139), .B(n2960), .Y(n3014) );
  CLKAND2X6 U108 ( .A(n2139), .B(n2961), .Y(n3016) );
  CLKAND2X6 U109 ( .A(n2139), .B(n2962), .Y(n3018) );
  CLKAND2X6 U110 ( .A(n2139), .B(n2963), .Y(n3019) );
  CLKAND2X6 U111 ( .A(n2139), .B(n2964), .Y(n3020) );
  CLKAND2X6 U112 ( .A(n2139), .B(n2965), .Y(n3021) );
  CLKAND2X6 U113 ( .A(n2139), .B(n2968), .Y(n3022) );
  CLKAND2X6 U114 ( .A(n2139), .B(n2979), .Y(n3023) );
  CLKAND2X6 U115 ( .A(n2139), .B(n2990), .Y(n3024) );
  INVXL U116 ( .A(n3120), .Y(n2133) );
  INVX6 U117 ( .A(n2133), .Y(n2134) );
  AND4X6 U118 ( .A(Jump[0]), .B(N1140), .C(n3101), .D(M[0]), .Y(n3036) );
  INVXL U119 ( .A(n3118), .Y(n2135) );
  INVX6 U120 ( .A(n46), .Y(n2137) );
  INVX6 U121 ( .A(n47), .Y(n2138) );
  INVX12 U122 ( .A(n43), .Y(n2139) );
  INVX12 U123 ( .A(n45), .Y(n2140) );
  INVXL U124 ( .A(n2927), .Y(n2141) );
  INVX12 U125 ( .A(n2141), .Y(n2142) );
  INVXL U126 ( .A(n2929), .Y(n2143) );
  INVX12 U127 ( .A(n2143), .Y(n2144) );
  INVXL U128 ( .A(n2930), .Y(n2145) );
  INVX12 U129 ( .A(n2145), .Y(n2146) );
  INVXL U130 ( .A(n2931), .Y(n2147) );
  INVX12 U131 ( .A(n2147), .Y(n2148) );
  INVXL U132 ( .A(n2932), .Y(n2149) );
  INVX12 U133 ( .A(n2149), .Y(n2150) );
  INVXL U134 ( .A(n2933), .Y(n2151) );
  INVX12 U135 ( .A(n2151), .Y(n2152) );
  INVXL U136 ( .A(n2934), .Y(n2153) );
  INVX12 U137 ( .A(n2153), .Y(n2154) );
  INVXL U138 ( .A(n2935), .Y(n2155) );
  INVX12 U139 ( .A(n2155), .Y(n2156) );
  INVXL U140 ( .A(n2936), .Y(n2157) );
  INVX12 U141 ( .A(n2157), .Y(n2158) );
  INVXL U142 ( .A(n2937), .Y(n2159) );
  INVX12 U143 ( .A(n2159), .Y(n2160) );
  INVXL U144 ( .A(n2938), .Y(n2161) );
  INVX12 U145 ( .A(n2161), .Y(n2162) );
  INVXL U146 ( .A(n2939), .Y(n2163) );
  INVX12 U147 ( .A(n2163), .Y(n2164) );
  INVXL U148 ( .A(n2940), .Y(n2165) );
  INVX12 U149 ( .A(n2165), .Y(n2166) );
  INVXL U150 ( .A(n2941), .Y(n2167) );
  INVX12 U151 ( .A(n2167), .Y(n2168) );
  INVXL U152 ( .A(n2942), .Y(n2169) );
  INVX12 U153 ( .A(n2169), .Y(n2170) );
  INVXL U154 ( .A(n2943), .Y(n2171) );
  INVX12 U155 ( .A(n2171), .Y(n2172) );
  INVXL U156 ( .A(n2944), .Y(n2173) );
  INVX12 U157 ( .A(n2173), .Y(n2174) );
  INVXL U158 ( .A(n2945), .Y(n2175) );
  INVX12 U159 ( .A(n2175), .Y(n2176) );
  INVXL U160 ( .A(n2946), .Y(n2177) );
  INVX12 U161 ( .A(n2177), .Y(n2178) );
  INVXL U162 ( .A(n2947), .Y(n2179) );
  INVX12 U163 ( .A(n2179), .Y(n2180) );
  INVXL U164 ( .A(n2948), .Y(n2181) );
  INVX12 U165 ( .A(n2181), .Y(n2182) );
  INVXL U166 ( .A(n2949), .Y(n2183) );
  INVX12 U167 ( .A(n2183), .Y(n2184) );
  INVXL U168 ( .A(n2950), .Y(n2185) );
  INVX12 U169 ( .A(n2185), .Y(n2186) );
  INVXL U170 ( .A(n2951), .Y(n2187) );
  INVX12 U171 ( .A(n2187), .Y(n2188) );
  INVXL U172 ( .A(n2952), .Y(n2189) );
  INVX12 U173 ( .A(n2189), .Y(n2190) );
  INVXL U174 ( .A(n2953), .Y(n2191) );
  INVX12 U175 ( .A(n2191), .Y(n2192) );
  INVXL U176 ( .A(n2954), .Y(n2193) );
  INVX12 U177 ( .A(n2193), .Y(n2194) );
  INVXL U178 ( .A(n2955), .Y(n2195) );
  INVX12 U179 ( .A(n2195), .Y(n2196) );
  INVXL U180 ( .A(n2956), .Y(n2197) );
  INVX12 U181 ( .A(n2197), .Y(n2198) );
  INVXL U182 ( .A(n2957), .Y(n2199) );
  INVX12 U183 ( .A(n2199), .Y(n2200) );
  INVXL U184 ( .A(n2958), .Y(n2201) );
  INVX12 U185 ( .A(n2201), .Y(n2202) );
  INVXL U186 ( .A(n2959), .Y(n2203) );
  INVX12 U187 ( .A(n2203), .Y(n2204) );
  CLKAND2X6 U188 ( .A(n3103), .B(n3004), .Y(n2966) );
  NOR3X2 U189 ( .A(n3110), .B(n3109), .C(n3107), .Y(n3004) );
  CLKAND2X6 U190 ( .A(n2993), .B(n2996), .Y(n2980) );
  NOR3X2 U191 ( .A(n3109), .B(WB_Rd[2]), .C(n3110), .Y(n2996) );
  CLKAND2X6 U192 ( .A(n3103), .B(n2996), .Y(n2971) );
  CLKAND2X6 U193 ( .A(n2993), .B(n3004), .Y(n2975) );
  CLKAND2X6 U194 ( .A(n3004), .B(n3005), .Y(n2984) );
  CLKAND2X6 U195 ( .A(n2996), .B(n3017), .Y(n2965) );
  CLKAND2X6 U196 ( .A(n2993), .B(n2998), .Y(n2981) );
  NOR3X2 U197 ( .A(WB_Rd[0]), .B(WB_Rd[2]), .C(n3110), .Y(n2998) );
  CLKAND2X6 U198 ( .A(n3103), .B(n3009), .Y(n2969) );
  NOR3X2 U199 ( .A(n3109), .B(WB_Rd[1]), .C(n3107), .Y(n3009) );
  CLKAND2X6 U200 ( .A(n2996), .B(n3005), .Y(n2988) );
  CLKAND2X6 U201 ( .A(n3004), .B(n3017), .Y(n2961) );
  CLKAND2X6 U202 ( .A(n2993), .B(n2994), .Y(n2978) );
  NOR3X2 U203 ( .A(WB_Rd[0]), .B(WB_Rd[1]), .C(n3107), .Y(n2994) );
  CLKAND2X6 U204 ( .A(n3103), .B(n3000), .Y(n2973) );
  NOR3X2 U205 ( .A(WB_Rd[1]), .B(WB_Rd[2]), .C(n3109), .Y(n3000) );
  CLKAND2X6 U206 ( .A(n2998), .B(n3017), .Y(n2968) );
  CLKAND2X6 U207 ( .A(n3009), .B(n3005), .Y(n2986) );
  CLKAND2X6 U208 ( .A(n2993), .B(n3007), .Y(n2976) );
  NOR3X2 U209 ( .A(n3110), .B(WB_Rd[0]), .C(n3107), .Y(n3007) );
  CLKAND2X6 U210 ( .A(n3103), .B(n3002), .Y(n2974) );
  CLKAND2X6 U211 ( .A(n2998), .B(n3005), .Y(n2989) );
  CLKAND2X6 U212 ( .A(n3009), .B(n3017), .Y(n2963) );
  CLKAND2X6 U213 ( .A(n3103), .B(n3007), .Y(n2967) );
  CLKAND2X6 U214 ( .A(n2993), .B(n3002), .Y(n2983) );
  CLKAND2X6 U215 ( .A(n2994), .B(n3017), .Y(n2964) );
  CLKAND2X6 U216 ( .A(n3000), .B(n3005), .Y(n2928) );
  CLKBUFX6 U217 ( .A(n3188), .Y(n2205) );
  CLKINVX2 U218 ( .A(PCWrite), .Y(n3116) );
  CLKAND2X6 U219 ( .A(n3103), .B(n2994), .Y(n2970) );
  CLKAND2X6 U220 ( .A(n2993), .B(n3000), .Y(n2982) );
  CLKAND2X6 U221 ( .A(n3007), .B(n3017), .Y(n2962) );
  CLKAND2X6 U222 ( .A(n3002), .B(n3005), .Y(n2960) );
  CLKBUFX6 U223 ( .A(n3185), .Y(n2206) );
  CLKBUFX6 U224 ( .A(n3187), .Y(n2207) );
  CLKMX2X12 U225 ( .A(after_B_mux[3]), .B(EX_signextend[3]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[3]) );
  CLKMX2X12 U226 ( .A(after_B_mux[1]), .B(EX_signextend[1]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[1]) );
  CLKMX2X12 U227 ( .A(after_B_mux[0]), .B(EX_signextend[0]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[0]) );
  INVX3 U228 ( .A(EX_reg[4]), .Y(n3026) );
  CLKAND2X6 U229 ( .A(n2993), .B(n3009), .Y(n2977) );
  CLKAND2X6 U230 ( .A(n2998), .B(n3103), .Y(n2972) );
  CLKAND2X6 U231 ( .A(n2994), .B(n3005), .Y(n2987) );
  CLKAND2X6 U232 ( .A(n3007), .B(n3005), .Y(n2985) );
  NOR3BX2 U233 ( .AN(WB_WB[0]), .B(n3015), .C(WB_Rd[4]), .Y(n3005) );
  CLKAND2X6 U234 ( .A(n3017), .B(n3000), .Y(n2979) );
  CLKAND2X6 U235 ( .A(n3017), .B(n3002), .Y(n2990) );
  NOR3BX2 U236 ( .AN(WB_WB[0]), .B(WB_Rd[3]), .C(WB_Rd[4]), .Y(n3017) );
  CLKBUFX6 U237 ( .A(n3183), .Y(n2208) );
  NOR2X6 U238 ( .A(WB_WB[1]), .B(WB_WB[2]), .Y(n3186) );
  CLKMX2X12 U239 ( .A(after_B_mux[5]), .B(EX_signextend[5]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[5]) );
  CLKMX2X12 U240 ( .A(after_B_mux[4]), .B(EX_signextend[4]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[4]) );
  CLKMX2X12 U241 ( .A(after_B_mux[2]), .B(EX_signextend[2]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[2]) );
  NOR2BXL U242 ( .AN(RegDST[0]), .B(n3116), .Y(EX_after_detect[4]) );
  INVXL U243 ( .A(DCACHE_addr[0]), .Y(n3137) );
  INVXL U244 ( .A(DCACHE_addr[1]), .Y(n3131) );
  INVXL U245 ( .A(DCACHE_addr[25]), .Y(n3143) );
  INVXL U246 ( .A(DCACHE_addr[24]), .Y(n3145) );
  INVXL U247 ( .A(DCACHE_addr[5]), .Y(n3123) );
  INVXL U248 ( .A(DCACHE_addr[6]), .Y(n3121) );
  INVXL U249 ( .A(DCACHE_addr[23]), .Y(n3147) );
  INVXL U250 ( .A(DCACHE_addr[7]), .Y(n3117) );
  INVXL U251 ( .A(DCACHE_addr[12]), .Y(n3171) );
  INVXL U252 ( .A(DCACHE_addr[17]), .Y(n3161) );
  INVXL U253 ( .A(DCACHE_addr[18]), .Y(n3157) );
  INVXL U254 ( .A(DCACHE_addr[19]), .Y(n3155) );
  INVXL U255 ( .A(DCACHE_addr[11]), .Y(n3173) );
  INVXL U256 ( .A(DCACHE_addr[13]), .Y(n3169) );
  INVXL U257 ( .A(DCACHE_addr[26]), .Y(n3141) );
  INVXL U258 ( .A(DCACHE_addr[29]), .Y(n3133) );
  INVXL U259 ( .A(DCACHE_addr[28]), .Y(n3135) );
  INVXL U260 ( .A(DCACHE_addr[9]), .Y(n3177) );
  INVXL U261 ( .A(DCACHE_addr[8]), .Y(n3179) );
  INVXL U262 ( .A(DCACHE_addr[21]), .Y(n3151) );
  INVXL U263 ( .A(DCACHE_addr[27]), .Y(n3139) );
  INVXL U264 ( .A(DCACHE_addr[15]), .Y(n3165) );
  INVXL U265 ( .A(DCACHE_addr[20]), .Y(n3153) );
  INVXL U266 ( .A(DCACHE_addr[22]), .Y(n3149) );
  INVXL U267 ( .A(DCACHE_addr[16]), .Y(n3163) );
  INVXL U268 ( .A(DCACHE_addr[10]), .Y(n3175) );
  INVXL U269 ( .A(DCACHE_addr[14]), .Y(n3167) );
  MXI4X1 U270 ( .A(\reg_file_next[24][6] ), .B(\reg_file_next[25][6] ), .C(
        \reg_file_next[26][6] ), .D(\reg_file_next[27][6] ), .S0(n2236), .S1(
        n2219), .Y(n2720) );
  MXI4X1 U271 ( .A(\reg_file_next[24][28] ), .B(\reg_file_next[25][28] ), .C(
        \reg_file_next[26][28] ), .D(\reg_file_next[27][28] ), .S0(n2231), 
        .S1(n2215), .Y(n2896) );
  MXI4X1 U272 ( .A(\reg_file_next[24][29] ), .B(\reg_file_next[25][29] ), .C(
        \reg_file_next[26][29] ), .D(\reg_file_next[27][29] ), .S0(n2231), 
        .S1(n2215), .Y(n2904) );
  MXI4X1 U273 ( .A(\reg_file_next[24][30] ), .B(\reg_file_next[25][30] ), .C(
        \reg_file_next[26][30] ), .D(\reg_file_next[27][30] ), .S0(n2232), 
        .S1(n2215), .Y(n2912) );
  MXI4X1 U274 ( .A(\reg_file_next[24][31] ), .B(\reg_file_next[25][31] ), .C(
        \reg_file_next[26][31] ), .D(\reg_file_next[27][31] ), .S0(n2232), 
        .S1(n2216), .Y(n2920) );
  MXI4X1 U275 ( .A(\reg_file_next[24][7] ), .B(\reg_file_next[25][7] ), .C(
        \reg_file_next[26][7] ), .D(\reg_file_next[27][7] ), .S0(n2237), .S1(
        n2219), .Y(n2728) );
  MXI4X1 U276 ( .A(\reg_file_next[24][8] ), .B(\reg_file_next[25][8] ), .C(
        \reg_file_next[26][8] ), .D(\reg_file_next[27][8] ), .S0(n2238), .S1(
        n2219), .Y(n2736) );
  MXI4X1 U277 ( .A(\reg_file_next[24][9] ), .B(\reg_file_next[25][9] ), .C(
        \reg_file_next[26][9] ), .D(\reg_file_next[27][9] ), .S0(n2238), .S1(
        n2220), .Y(n2744) );
  MXI4X1 U278 ( .A(\reg_file_next[24][10] ), .B(\reg_file_next[25][10] ), .C(
        \reg_file_next[26][10] ), .D(\reg_file_next[27][10] ), .S0(n2239), 
        .S1(n2220), .Y(n2752) );
  MXI4X1 U279 ( .A(\reg_file_next[24][11] ), .B(\reg_file_next[25][11] ), .C(
        \reg_file_next[26][11] ), .D(\reg_file_next[27][11] ), .S0(n2239), 
        .S1(n2221), .Y(n2760) );
  MXI4X1 U280 ( .A(\reg_file_next[24][12] ), .B(\reg_file_next[25][12] ), .C(
        \reg_file_next[26][12] ), .D(\reg_file_next[27][12] ), .S0(n2240), 
        .S1(n2221), .Y(n2768) );
  MXI4X1 U281 ( .A(\reg_file_next[24][13] ), .B(\reg_file_next[25][13] ), .C(
        \reg_file_next[26][13] ), .D(\reg_file_next[27][13] ), .S0(n2240), 
        .S1(n2221), .Y(n2776) );
  MXI4X1 U282 ( .A(\reg_file_next[24][14] ), .B(\reg_file_next[25][14] ), .C(
        \reg_file_next[26][14] ), .D(\reg_file_next[27][14] ), .S0(n2241), 
        .S1(n2222), .Y(n2784) );
  MXI4X1 U283 ( .A(\reg_file_next[24][15] ), .B(\reg_file_next[25][15] ), .C(
        \reg_file_next[26][15] ), .D(\reg_file_next[27][15] ), .S0(n2224), 
        .S1(n2222), .Y(n2792) );
  MXI4X1 U284 ( .A(\reg_file_next[24][16] ), .B(\reg_file_next[25][16] ), .C(
        \reg_file_next[26][16] ), .D(\reg_file_next[27][16] ), .S0(n2224), 
        .S1(n2210), .Y(n2800) );
  MXI4X1 U285 ( .A(\reg_file_next[24][17] ), .B(\reg_file_next[25][17] ), .C(
        \reg_file_next[26][17] ), .D(\reg_file_next[27][17] ), .S0(n2224), 
        .S1(n2210), .Y(n2808) );
  MXI4X1 U286 ( .A(\reg_file_next[24][18] ), .B(\reg_file_next[25][18] ), .C(
        \reg_file_next[26][18] ), .D(\reg_file_next[27][18] ), .S0(n2225), 
        .S1(n2211), .Y(n2816) );
  MXI4X1 U287 ( .A(\reg_file_next[24][19] ), .B(\reg_file_next[25][19] ), .C(
        \reg_file_next[26][19] ), .D(\reg_file_next[27][19] ), .S0(n2226), 
        .S1(n2211), .Y(n2824) );
  MXI4X1 U288 ( .A(\reg_file_next[24][20] ), .B(\reg_file_next[25][20] ), .C(
        \reg_file_next[26][20] ), .D(\reg_file_next[27][20] ), .S0(n2226), 
        .S1(n2211), .Y(n2832) );
  MXI4X1 U289 ( .A(\reg_file_next[24][21] ), .B(\reg_file_next[25][21] ), .C(
        \reg_file_next[26][21] ), .D(\reg_file_next[27][21] ), .S0(n2227), 
        .S1(n2212), .Y(n2840) );
  MXI4X1 U290 ( .A(\reg_file_next[24][22] ), .B(\reg_file_next[25][22] ), .C(
        \reg_file_next[26][22] ), .D(\reg_file_next[27][22] ), .S0(n2227), 
        .S1(n2212), .Y(n2848) );
  MXI4X1 U291 ( .A(\reg_file_next[24][23] ), .B(\reg_file_next[25][23] ), .C(
        \reg_file_next[26][23] ), .D(\reg_file_next[27][23] ), .S0(n2228), 
        .S1(n2213), .Y(n2856) );
  MXI4X1 U292 ( .A(\reg_file_next[24][24] ), .B(\reg_file_next[25][24] ), .C(
        \reg_file_next[26][24] ), .D(\reg_file_next[27][24] ), .S0(n2228), 
        .S1(n2213), .Y(n2864) );
  MXI4X1 U293 ( .A(\reg_file_next[24][25] ), .B(\reg_file_next[25][25] ), .C(
        \reg_file_next[26][25] ), .D(\reg_file_next[27][25] ), .S0(n2229), 
        .S1(n2213), .Y(n2872) );
  MXI4X1 U294 ( .A(\reg_file_next[24][26] ), .B(\reg_file_next[25][26] ), .C(
        \reg_file_next[26][26] ), .D(\reg_file_next[27][26] ), .S0(n2230), 
        .S1(n2214), .Y(n2880) );
  MXI4X1 U295 ( .A(\reg_file_next[24][27] ), .B(\reg_file_next[25][27] ), .C(
        \reg_file_next[26][27] ), .D(\reg_file_next[27][27] ), .S0(n2230), 
        .S1(n2214), .Y(n2888) );
  NOR2BXL U296 ( .AN(\MemtoReg[0] ), .B(n3116), .Y(WB_after_detect[1]) );
  MXI2XL U297 ( .A(n1874), .B(n2204), .S0(n2961), .Y(\reg_file_next[7][0] ) );
  MXI2XL U298 ( .A(n2002), .B(n2204), .S0(n2965), .Y(\reg_file_next[3][0] ) );
  MXI2XL U299 ( .A(n1618), .B(n2204), .S0(n2984), .Y(\reg_file_next[15][0] )
         );
  MXI2XL U300 ( .A(n1746), .B(n2204), .S0(n2988), .Y(\reg_file_next[11][0] )
         );
  MXI2XL U301 ( .A(n1362), .B(n2204), .S0(n2975), .Y(\reg_file_next[23][0] )
         );
  MXI2XL U302 ( .A(n1490), .B(n2204), .S0(n2980), .Y(\reg_file_next[19][0] )
         );
  MXI2XL U303 ( .A(n49), .B(n2204), .S0(n2966), .Y(\reg_file_next[31][0] ) );
  MXI2XL U304 ( .A(n1875), .B(n2182), .S0(n2961), .Y(\reg_file_next[7][1] ) );
  MXI2XL U305 ( .A(n2003), .B(n2182), .S0(n2965), .Y(\reg_file_next[3][1] ) );
  MXI2XL U306 ( .A(n1619), .B(n2182), .S0(n2984), .Y(\reg_file_next[15][1] )
         );
  MXI2XL U307 ( .A(n1747), .B(n2182), .S0(n2988), .Y(\reg_file_next[11][1] )
         );
  MXI2XL U308 ( .A(n1363), .B(n2182), .S0(n2975), .Y(\reg_file_next[23][1] )
         );
  MXI2XL U309 ( .A(n1491), .B(n2182), .S0(n2980), .Y(\reg_file_next[19][1] )
         );
  MXI2XL U310 ( .A(n50), .B(n2182), .S0(n2966), .Y(\reg_file_next[31][1] ) );
  MXI2XL U311 ( .A(n1876), .B(n2160), .S0(n2961), .Y(\reg_file_next[7][2] ) );
  MXI2XL U312 ( .A(n2004), .B(n2160), .S0(n2965), .Y(\reg_file_next[3][2] ) );
  MXI2XL U313 ( .A(n1620), .B(n2160), .S0(n2984), .Y(\reg_file_next[15][2] )
         );
  MXI2XL U314 ( .A(n1748), .B(n2160), .S0(n2988), .Y(\reg_file_next[11][2] )
         );
  MXI2XL U315 ( .A(n1364), .B(n2160), .S0(n2975), .Y(\reg_file_next[23][2] )
         );
  MXI2XL U316 ( .A(n1492), .B(n2160), .S0(n2980), .Y(\reg_file_next[19][2] )
         );
  MXI2XL U317 ( .A(n51), .B(n2160), .S0(n2966), .Y(\reg_file_next[31][2] ) );
  MXI2XL U318 ( .A(n1877), .B(n2154), .S0(n2961), .Y(\reg_file_next[7][3] ) );
  MXI2XL U319 ( .A(n2005), .B(n2154), .S0(n2965), .Y(\reg_file_next[3][3] ) );
  MXI2XL U320 ( .A(n1621), .B(n2154), .S0(n2984), .Y(\reg_file_next[15][3] )
         );
  MXI2XL U321 ( .A(n1749), .B(n2154), .S0(n2988), .Y(\reg_file_next[11][3] )
         );
  MXI2XL U322 ( .A(n1365), .B(n2154), .S0(n2975), .Y(\reg_file_next[23][3] )
         );
  MXI2XL U323 ( .A(n1493), .B(n2154), .S0(n2980), .Y(\reg_file_next[19][3] )
         );
  MXI2XL U324 ( .A(n52), .B(n2154), .S0(n2966), .Y(\reg_file_next[31][3] ) );
  MXI2XL U325 ( .A(n1878), .B(n2152), .S0(n2961), .Y(\reg_file_next[7][4] ) );
  MXI2XL U326 ( .A(n2006), .B(n2152), .S0(n2965), .Y(\reg_file_next[3][4] ) );
  MXI2XL U327 ( .A(n1622), .B(n2152), .S0(n2984), .Y(\reg_file_next[15][4] )
         );
  MXI2XL U328 ( .A(n1750), .B(n2152), .S0(n2988), .Y(\reg_file_next[11][4] )
         );
  MXI2XL U329 ( .A(n1366), .B(n2152), .S0(n2975), .Y(\reg_file_next[23][4] )
         );
  MXI2XL U330 ( .A(n1494), .B(n2152), .S0(n2980), .Y(\reg_file_next[19][4] )
         );
  MXI2XL U331 ( .A(n53), .B(n2152), .S0(n2966), .Y(\reg_file_next[31][4] ) );
  MXI2XL U332 ( .A(n1879), .B(n2150), .S0(n2961), .Y(\reg_file_next[7][5] ) );
  MXI2XL U333 ( .A(n2007), .B(n2150), .S0(n2965), .Y(\reg_file_next[3][5] ) );
  MXI2XL U334 ( .A(n1623), .B(n2150), .S0(n2984), .Y(\reg_file_next[15][5] )
         );
  MXI2XL U335 ( .A(n1751), .B(n2150), .S0(n2988), .Y(\reg_file_next[11][5] )
         );
  MXI2XL U336 ( .A(n1367), .B(n2150), .S0(n2975), .Y(\reg_file_next[23][5] )
         );
  MXI2XL U337 ( .A(n1495), .B(n2150), .S0(n2980), .Y(\reg_file_next[19][5] )
         );
  MXI2XL U338 ( .A(n54), .B(n2150), .S0(n2966), .Y(\reg_file_next[31][5] ) );
  MXI2XL U339 ( .A(n1880), .B(n2148), .S0(n2961), .Y(\reg_file_next[7][6] ) );
  MXI2XL U340 ( .A(n2008), .B(n2148), .S0(n2965), .Y(\reg_file_next[3][6] ) );
  MXI2XL U341 ( .A(n1624), .B(n2148), .S0(n2984), .Y(\reg_file_next[15][6] )
         );
  MXI2XL U342 ( .A(n1752), .B(n2148), .S0(n2988), .Y(\reg_file_next[11][6] )
         );
  MXI2XL U343 ( .A(n1368), .B(n2148), .S0(n2975), .Y(\reg_file_next[23][6] )
         );
  MXI2XL U344 ( .A(n1496), .B(n2148), .S0(n2980), .Y(\reg_file_next[19][6] )
         );
  MXI2XL U345 ( .A(n55), .B(n2148), .S0(n2966), .Y(\reg_file_next[31][6] ) );
  MXI2XL U346 ( .A(n1881), .B(n2146), .S0(n2961), .Y(\reg_file_next[7][7] ) );
  MXI2XL U347 ( .A(n2009), .B(n2146), .S0(n2965), .Y(\reg_file_next[3][7] ) );
  MXI2XL U348 ( .A(n1625), .B(n2146), .S0(n2984), .Y(\reg_file_next[15][7] )
         );
  MXI2XL U349 ( .A(n1753), .B(n2146), .S0(n2988), .Y(\reg_file_next[11][7] )
         );
  MXI2XL U350 ( .A(n1369), .B(n2146), .S0(n2975), .Y(\reg_file_next[23][7] )
         );
  MXI2XL U351 ( .A(n1497), .B(n2146), .S0(n2980), .Y(\reg_file_next[19][7] )
         );
  MXI2XL U352 ( .A(n56), .B(n2146), .S0(n2966), .Y(\reg_file_next[31][7] ) );
  MXI2XL U353 ( .A(n1882), .B(n2144), .S0(n2961), .Y(\reg_file_next[7][8] ) );
  MXI2XL U354 ( .A(n2010), .B(n2144), .S0(n2965), .Y(\reg_file_next[3][8] ) );
  MXI2XL U355 ( .A(n1626), .B(n2144), .S0(n2984), .Y(\reg_file_next[15][8] )
         );
  MXI2XL U356 ( .A(n1754), .B(n2144), .S0(n2988), .Y(\reg_file_next[11][8] )
         );
  MXI2XL U357 ( .A(n1370), .B(n2144), .S0(n2975), .Y(\reg_file_next[23][8] )
         );
  MXI2XL U358 ( .A(n1498), .B(n2144), .S0(n2980), .Y(\reg_file_next[19][8] )
         );
  MXI2XL U359 ( .A(n57), .B(n2144), .S0(n2966), .Y(\reg_file_next[31][8] ) );
  MXI2XL U360 ( .A(n1883), .B(n2142), .S0(n2961), .Y(\reg_file_next[7][9] ) );
  MXI2XL U361 ( .A(n2011), .B(n2142), .S0(n2965), .Y(\reg_file_next[3][9] ) );
  MXI2XL U362 ( .A(n1627), .B(n2142), .S0(n2984), .Y(\reg_file_next[15][9] )
         );
  MXI2XL U363 ( .A(n1755), .B(n2142), .S0(n2988), .Y(\reg_file_next[11][9] )
         );
  MXI2XL U364 ( .A(n1371), .B(n2142), .S0(n2975), .Y(\reg_file_next[23][9] )
         );
  MXI2XL U365 ( .A(n1499), .B(n2142), .S0(n2980), .Y(\reg_file_next[19][9] )
         );
  MXI2XL U366 ( .A(n58), .B(n2142), .S0(n2966), .Y(\reg_file_next[31][9] ) );
  MXI2XL U367 ( .A(n1884), .B(n2202), .S0(n2961), .Y(\reg_file_next[7][10] )
         );
  MXI2XL U368 ( .A(n2012), .B(n2202), .S0(n2965), .Y(\reg_file_next[3][10] )
         );
  MXI2XL U369 ( .A(n1628), .B(n2202), .S0(n2984), .Y(\reg_file_next[15][10] )
         );
  MXI2XL U370 ( .A(n1756), .B(n2202), .S0(n2988), .Y(\reg_file_next[11][10] )
         );
  MXI2XL U371 ( .A(n1372), .B(n2202), .S0(n2975), .Y(\reg_file_next[23][10] )
         );
  MXI2XL U372 ( .A(n1500), .B(n2202), .S0(n2980), .Y(\reg_file_next[19][10] )
         );
  MXI2XL U373 ( .A(n59), .B(n2202), .S0(n2966), .Y(\reg_file_next[31][10] ) );
  MXI2XL U374 ( .A(n1885), .B(n2200), .S0(n2961), .Y(\reg_file_next[7][11] )
         );
  MXI2XL U375 ( .A(n2013), .B(n2200), .S0(n2965), .Y(\reg_file_next[3][11] )
         );
  MXI2XL U376 ( .A(n1629), .B(n2200), .S0(n2984), .Y(\reg_file_next[15][11] )
         );
  MXI2XL U377 ( .A(n1757), .B(n2200), .S0(n2988), .Y(\reg_file_next[11][11] )
         );
  MXI2XL U378 ( .A(n1373), .B(n2200), .S0(n2975), .Y(\reg_file_next[23][11] )
         );
  MXI2XL U379 ( .A(n1501), .B(n2200), .S0(n2980), .Y(\reg_file_next[19][11] )
         );
  MXI2XL U380 ( .A(n60), .B(n2200), .S0(n2966), .Y(\reg_file_next[31][11] ) );
  MXI2XL U381 ( .A(n1886), .B(n2198), .S0(n2961), .Y(\reg_file_next[7][12] )
         );
  MXI2XL U382 ( .A(n2014), .B(n2198), .S0(n2965), .Y(\reg_file_next[3][12] )
         );
  MXI2XL U383 ( .A(n1630), .B(n2198), .S0(n2984), .Y(\reg_file_next[15][12] )
         );
  MXI2XL U384 ( .A(n1758), .B(n2198), .S0(n2988), .Y(\reg_file_next[11][12] )
         );
  MXI2XL U385 ( .A(n1374), .B(n2198), .S0(n2975), .Y(\reg_file_next[23][12] )
         );
  MXI2XL U386 ( .A(n1502), .B(n2198), .S0(n2980), .Y(\reg_file_next[19][12] )
         );
  MXI2XL U387 ( .A(n61), .B(n2198), .S0(n2966), .Y(\reg_file_next[31][12] ) );
  MXI2XL U388 ( .A(n1887), .B(n2196), .S0(n2961), .Y(\reg_file_next[7][13] )
         );
  MXI2XL U389 ( .A(n2015), .B(n2196), .S0(n2965), .Y(\reg_file_next[3][13] )
         );
  MXI2XL U390 ( .A(n1631), .B(n2196), .S0(n2984), .Y(\reg_file_next[15][13] )
         );
  MXI2XL U391 ( .A(n1759), .B(n2196), .S0(n2988), .Y(\reg_file_next[11][13] )
         );
  MXI2XL U392 ( .A(n1375), .B(n2196), .S0(n2975), .Y(\reg_file_next[23][13] )
         );
  MXI2XL U393 ( .A(n1503), .B(n2196), .S0(n2980), .Y(\reg_file_next[19][13] )
         );
  MXI2XL U394 ( .A(n62), .B(n2196), .S0(n2966), .Y(\reg_file_next[31][13] ) );
  MXI2XL U395 ( .A(n1888), .B(n2194), .S0(n2961), .Y(\reg_file_next[7][14] )
         );
  MXI2XL U396 ( .A(n2016), .B(n2194), .S0(n2965), .Y(\reg_file_next[3][14] )
         );
  MXI2XL U397 ( .A(n1632), .B(n2194), .S0(n2984), .Y(\reg_file_next[15][14] )
         );
  MXI2XL U398 ( .A(n1760), .B(n2194), .S0(n2988), .Y(\reg_file_next[11][14] )
         );
  MXI2XL U399 ( .A(n1376), .B(n2194), .S0(n2975), .Y(\reg_file_next[23][14] )
         );
  MXI2XL U400 ( .A(n1504), .B(n2194), .S0(n2980), .Y(\reg_file_next[19][14] )
         );
  MXI2XL U401 ( .A(n63), .B(n2194), .S0(n2966), .Y(\reg_file_next[31][14] ) );
  MXI2XL U402 ( .A(n1889), .B(n2192), .S0(n2961), .Y(\reg_file_next[7][15] )
         );
  MXI2XL U403 ( .A(n2017), .B(n2192), .S0(n2965), .Y(\reg_file_next[3][15] )
         );
  MXI2XL U404 ( .A(n1633), .B(n2192), .S0(n2984), .Y(\reg_file_next[15][15] )
         );
  MXI2XL U405 ( .A(n1761), .B(n2192), .S0(n2988), .Y(\reg_file_next[11][15] )
         );
  MXI2XL U406 ( .A(n1377), .B(n2192), .S0(n2975), .Y(\reg_file_next[23][15] )
         );
  MXI2XL U407 ( .A(n1505), .B(n2192), .S0(n2980), .Y(\reg_file_next[19][15] )
         );
  MXI2XL U408 ( .A(n64), .B(n2192), .S0(n2966), .Y(\reg_file_next[31][15] ) );
  MXI2XL U409 ( .A(n1890), .B(n2190), .S0(n2961), .Y(\reg_file_next[7][16] )
         );
  MXI2XL U410 ( .A(n2018), .B(n2190), .S0(n2965), .Y(\reg_file_next[3][16] )
         );
  MXI2XL U411 ( .A(n1634), .B(n2190), .S0(n2984), .Y(\reg_file_next[15][16] )
         );
  MXI2XL U412 ( .A(n1762), .B(n2190), .S0(n2988), .Y(\reg_file_next[11][16] )
         );
  MXI2XL U413 ( .A(n1378), .B(n2190), .S0(n2975), .Y(\reg_file_next[23][16] )
         );
  MXI2XL U414 ( .A(n1506), .B(n2190), .S0(n2980), .Y(\reg_file_next[19][16] )
         );
  MXI2XL U415 ( .A(n65), .B(n2190), .S0(n2966), .Y(\reg_file_next[31][16] ) );
  MXI2XL U416 ( .A(n1891), .B(n2188), .S0(n2961), .Y(\reg_file_next[7][17] )
         );
  MXI2XL U417 ( .A(n2019), .B(n2188), .S0(n2965), .Y(\reg_file_next[3][17] )
         );
  MXI2XL U418 ( .A(n1635), .B(n2188), .S0(n2984), .Y(\reg_file_next[15][17] )
         );
  MXI2XL U419 ( .A(n1763), .B(n2188), .S0(n2988), .Y(\reg_file_next[11][17] )
         );
  MXI2XL U420 ( .A(n1379), .B(n2188), .S0(n2975), .Y(\reg_file_next[23][17] )
         );
  MXI2XL U421 ( .A(n1507), .B(n2188), .S0(n2980), .Y(\reg_file_next[19][17] )
         );
  MXI2XL U422 ( .A(n66), .B(n2188), .S0(n2966), .Y(\reg_file_next[31][17] ) );
  MXI2XL U423 ( .A(n1892), .B(n2186), .S0(n2961), .Y(\reg_file_next[7][18] )
         );
  MXI2XL U424 ( .A(n2020), .B(n2186), .S0(n2965), .Y(\reg_file_next[3][18] )
         );
  MXI2XL U425 ( .A(n1636), .B(n2186), .S0(n2984), .Y(\reg_file_next[15][18] )
         );
  MXI2XL U426 ( .A(n1764), .B(n2186), .S0(n2988), .Y(\reg_file_next[11][18] )
         );
  MXI2XL U427 ( .A(n1380), .B(n2186), .S0(n2975), .Y(\reg_file_next[23][18] )
         );
  MXI2XL U428 ( .A(n1508), .B(n2186), .S0(n2980), .Y(\reg_file_next[19][18] )
         );
  MXI2XL U429 ( .A(n67), .B(n2186), .S0(n2966), .Y(\reg_file_next[31][18] ) );
  MXI2XL U430 ( .A(n1893), .B(n2184), .S0(n2961), .Y(\reg_file_next[7][19] )
         );
  MXI2XL U431 ( .A(n2021), .B(n2184), .S0(n2965), .Y(\reg_file_next[3][19] )
         );
  MXI2XL U432 ( .A(n1637), .B(n2184), .S0(n2984), .Y(\reg_file_next[15][19] )
         );
  MXI2XL U433 ( .A(n1765), .B(n2184), .S0(n2988), .Y(\reg_file_next[11][19] )
         );
  MXI2XL U434 ( .A(n1381), .B(n2184), .S0(n2975), .Y(\reg_file_next[23][19] )
         );
  MXI2XL U435 ( .A(n1509), .B(n2184), .S0(n2980), .Y(\reg_file_next[19][19] )
         );
  MXI2XL U436 ( .A(n68), .B(n2184), .S0(n2966), .Y(\reg_file_next[31][19] ) );
  MXI2XL U437 ( .A(n1894), .B(n2180), .S0(n2961), .Y(\reg_file_next[7][20] )
         );
  MXI2XL U438 ( .A(n2022), .B(n2180), .S0(n2965), .Y(\reg_file_next[3][20] )
         );
  MXI2XL U439 ( .A(n1638), .B(n2180), .S0(n2984), .Y(\reg_file_next[15][20] )
         );
  MXI2XL U440 ( .A(n1766), .B(n2180), .S0(n2988), .Y(\reg_file_next[11][20] )
         );
  MXI2XL U441 ( .A(n1382), .B(n2180), .S0(n2975), .Y(\reg_file_next[23][20] )
         );
  MXI2XL U442 ( .A(n1510), .B(n2180), .S0(n2980), .Y(\reg_file_next[19][20] )
         );
  MXI2XL U443 ( .A(n69), .B(n2180), .S0(n2966), .Y(\reg_file_next[31][20] ) );
  MXI2XL U444 ( .A(n1895), .B(n2178), .S0(n2961), .Y(\reg_file_next[7][21] )
         );
  MXI2XL U445 ( .A(n2023), .B(n2178), .S0(n2965), .Y(\reg_file_next[3][21] )
         );
  MXI2XL U446 ( .A(n1639), .B(n2178), .S0(n2984), .Y(\reg_file_next[15][21] )
         );
  MXI2XL U447 ( .A(n1767), .B(n2178), .S0(n2988), .Y(\reg_file_next[11][21] )
         );
  MXI2XL U448 ( .A(n1383), .B(n2178), .S0(n2975), .Y(\reg_file_next[23][21] )
         );
  MXI2XL U449 ( .A(n1511), .B(n2178), .S0(n2980), .Y(\reg_file_next[19][21] )
         );
  MXI2XL U450 ( .A(n71), .B(n2178), .S0(n2966), .Y(\reg_file_next[31][21] ) );
  MXI2XL U451 ( .A(n1896), .B(n2176), .S0(n2961), .Y(\reg_file_next[7][22] )
         );
  MXI2XL U452 ( .A(n2024), .B(n2176), .S0(n2965), .Y(\reg_file_next[3][22] )
         );
  MXI2XL U453 ( .A(n1640), .B(n2176), .S0(n2984), .Y(\reg_file_next[15][22] )
         );
  MXI2XL U454 ( .A(n1768), .B(n2176), .S0(n2988), .Y(\reg_file_next[11][22] )
         );
  MXI2XL U455 ( .A(n1384), .B(n2176), .S0(n2975), .Y(\reg_file_next[23][22] )
         );
  MXI2XL U456 ( .A(n1512), .B(n2176), .S0(n2980), .Y(\reg_file_next[19][22] )
         );
  MXI2XL U457 ( .A(n72), .B(n2176), .S0(n2966), .Y(\reg_file_next[31][22] ) );
  MXI2XL U458 ( .A(n1897), .B(n2174), .S0(n2961), .Y(\reg_file_next[7][23] )
         );
  MXI2XL U459 ( .A(n2025), .B(n2174), .S0(n2965), .Y(\reg_file_next[3][23] )
         );
  MXI2XL U460 ( .A(n1641), .B(n2174), .S0(n2984), .Y(\reg_file_next[15][23] )
         );
  MXI2XL U461 ( .A(n1769), .B(n2174), .S0(n2988), .Y(\reg_file_next[11][23] )
         );
  MXI2XL U462 ( .A(n1385), .B(n2174), .S0(n2975), .Y(\reg_file_next[23][23] )
         );
  MXI2XL U463 ( .A(n1513), .B(n2174), .S0(n2980), .Y(\reg_file_next[19][23] )
         );
  MXI2XL U464 ( .A(n73), .B(n2174), .S0(n2966), .Y(\reg_file_next[31][23] ) );
  MXI2XL U465 ( .A(n1898), .B(n2172), .S0(n2961), .Y(\reg_file_next[7][24] )
         );
  MXI2XL U466 ( .A(n2026), .B(n2172), .S0(n2965), .Y(\reg_file_next[3][24] )
         );
  MXI2XL U467 ( .A(n1642), .B(n2172), .S0(n2984), .Y(\reg_file_next[15][24] )
         );
  MXI2XL U468 ( .A(n1770), .B(n2172), .S0(n2988), .Y(\reg_file_next[11][24] )
         );
  MXI2XL U469 ( .A(n1386), .B(n2172), .S0(n2975), .Y(\reg_file_next[23][24] )
         );
  MXI2XL U470 ( .A(n1514), .B(n2172), .S0(n2980), .Y(\reg_file_next[19][24] )
         );
  MXI2XL U471 ( .A(n74), .B(n2172), .S0(n2966), .Y(\reg_file_next[31][24] ) );
  MXI2XL U472 ( .A(n1899), .B(n2170), .S0(n2961), .Y(\reg_file_next[7][25] )
         );
  MXI2XL U473 ( .A(n2027), .B(n2170), .S0(n2965), .Y(\reg_file_next[3][25] )
         );
  MXI2XL U474 ( .A(n1643), .B(n2170), .S0(n2984), .Y(\reg_file_next[15][25] )
         );
  MXI2XL U475 ( .A(n1771), .B(n2170), .S0(n2988), .Y(\reg_file_next[11][25] )
         );
  MXI2XL U476 ( .A(n1387), .B(n2170), .S0(n2975), .Y(\reg_file_next[23][25] )
         );
  MXI2XL U477 ( .A(n1515), .B(n2170), .S0(n2980), .Y(\reg_file_next[19][25] )
         );
  MXI2XL U478 ( .A(n75), .B(n2170), .S0(n2966), .Y(\reg_file_next[31][25] ) );
  MXI2XL U479 ( .A(n1900), .B(n2168), .S0(n2961), .Y(\reg_file_next[7][26] )
         );
  MXI2XL U480 ( .A(n2028), .B(n2168), .S0(n2965), .Y(\reg_file_next[3][26] )
         );
  MXI2XL U481 ( .A(n1644), .B(n2168), .S0(n2984), .Y(\reg_file_next[15][26] )
         );
  MXI2XL U482 ( .A(n1772), .B(n2168), .S0(n2988), .Y(\reg_file_next[11][26] )
         );
  MXI2XL U483 ( .A(n1388), .B(n2168), .S0(n2975), .Y(\reg_file_next[23][26] )
         );
  MXI2XL U484 ( .A(n1516), .B(n2168), .S0(n2980), .Y(\reg_file_next[19][26] )
         );
  MXI2XL U485 ( .A(n76), .B(n2168), .S0(n2966), .Y(\reg_file_next[31][26] ) );
  MXI2XL U486 ( .A(n1901), .B(n2166), .S0(n2961), .Y(\reg_file_next[7][27] )
         );
  MXI2XL U487 ( .A(n2029), .B(n2166), .S0(n2965), .Y(\reg_file_next[3][27] )
         );
  MXI2XL U488 ( .A(n1645), .B(n2166), .S0(n2984), .Y(\reg_file_next[15][27] )
         );
  MXI2XL U489 ( .A(n1773), .B(n2166), .S0(n2988), .Y(\reg_file_next[11][27] )
         );
  MXI2XL U490 ( .A(n1389), .B(n2166), .S0(n2975), .Y(\reg_file_next[23][27] )
         );
  MXI2XL U491 ( .A(n1517), .B(n2166), .S0(n2980), .Y(\reg_file_next[19][27] )
         );
  MXI2XL U492 ( .A(n77), .B(n2166), .S0(n2966), .Y(\reg_file_next[31][27] ) );
  MXI2XL U493 ( .A(n1902), .B(n2164), .S0(n2961), .Y(\reg_file_next[7][28] )
         );
  MXI2XL U494 ( .A(n2030), .B(n2164), .S0(n2965), .Y(\reg_file_next[3][28] )
         );
  MXI2XL U495 ( .A(n1646), .B(n2164), .S0(n2984), .Y(\reg_file_next[15][28] )
         );
  MXI2XL U496 ( .A(n1774), .B(n2164), .S0(n2988), .Y(\reg_file_next[11][28] )
         );
  MXI2XL U497 ( .A(n1390), .B(n2164), .S0(n2975), .Y(\reg_file_next[23][28] )
         );
  MXI2XL U498 ( .A(n1518), .B(n2164), .S0(n2980), .Y(\reg_file_next[19][28] )
         );
  MXI2XL U499 ( .A(n78), .B(n2164), .S0(n2966), .Y(\reg_file_next[31][28] ) );
  MXI2XL U500 ( .A(n1903), .B(n2162), .S0(n2961), .Y(\reg_file_next[7][29] )
         );
  MXI2XL U501 ( .A(n2031), .B(n2162), .S0(n2965), .Y(\reg_file_next[3][29] )
         );
  MXI2XL U502 ( .A(n1647), .B(n2162), .S0(n2984), .Y(\reg_file_next[15][29] )
         );
  MXI2XL U503 ( .A(n1775), .B(n2162), .S0(n2988), .Y(\reg_file_next[11][29] )
         );
  MXI2XL U504 ( .A(n1391), .B(n2162), .S0(n2975), .Y(\reg_file_next[23][29] )
         );
  MXI2XL U505 ( .A(n1519), .B(n2162), .S0(n2980), .Y(\reg_file_next[19][29] )
         );
  MXI2XL U506 ( .A(n79), .B(n2162), .S0(n2966), .Y(\reg_file_next[31][29] ) );
  MXI2XL U507 ( .A(n1904), .B(n2158), .S0(n2961), .Y(\reg_file_next[7][30] )
         );
  MXI2XL U508 ( .A(n2032), .B(n2158), .S0(n2965), .Y(\reg_file_next[3][30] )
         );
  MXI2XL U509 ( .A(n1648), .B(n2158), .S0(n2984), .Y(\reg_file_next[15][30] )
         );
  MXI2XL U510 ( .A(n1776), .B(n2158), .S0(n2988), .Y(\reg_file_next[11][30] )
         );
  MXI2XL U511 ( .A(n1392), .B(n2158), .S0(n2975), .Y(\reg_file_next[23][30] )
         );
  MXI2XL U512 ( .A(n1520), .B(n2158), .S0(n2980), .Y(\reg_file_next[19][30] )
         );
  MXI2XL U513 ( .A(n80), .B(n2158), .S0(n2966), .Y(\reg_file_next[31][30] ) );
  MXI2XL U514 ( .A(n1905), .B(n2156), .S0(n2961), .Y(\reg_file_next[7][31] )
         );
  MXI2XL U515 ( .A(n2033), .B(n2156), .S0(n2965), .Y(\reg_file_next[3][31] )
         );
  MXI2XL U516 ( .A(n1649), .B(n2156), .S0(n2984), .Y(\reg_file_next[15][31] )
         );
  MXI2XL U517 ( .A(n1777), .B(n2156), .S0(n2988), .Y(\reg_file_next[11][31] )
         );
  MXI2XL U518 ( .A(n1393), .B(n2156), .S0(n2975), .Y(\reg_file_next[23][31] )
         );
  MXI2XL U519 ( .A(n1521), .B(n2156), .S0(n2980), .Y(\reg_file_next[19][31] )
         );
  MXI2XL U520 ( .A(n81), .B(n2156), .S0(n2966), .Y(\reg_file_next[31][31] ) );
  MXI2XL U521 ( .A(n178), .B(n2204), .S0(n2971), .Y(\reg_file_next[27][0] ) );
  MXI2XL U522 ( .A(n179), .B(n2182), .S0(n2971), .Y(\reg_file_next[27][1] ) );
  MXI2XL U523 ( .A(n180), .B(n2160), .S0(n2971), .Y(\reg_file_next[27][2] ) );
  MXI2XL U524 ( .A(n181), .B(n2154), .S0(n2971), .Y(\reg_file_next[27][3] ) );
  MXI2XL U525 ( .A(n182), .B(n2152), .S0(n2971), .Y(\reg_file_next[27][4] ) );
  MXI2XL U526 ( .A(n183), .B(n2150), .S0(n2971), .Y(\reg_file_next[27][5] ) );
  MXI2XL U527 ( .A(n184), .B(n2148), .S0(n2971), .Y(\reg_file_next[27][6] ) );
  MXI2XL U528 ( .A(n185), .B(n2146), .S0(n2971), .Y(\reg_file_next[27][7] ) );
  MXI2XL U529 ( .A(n186), .B(n2144), .S0(n2971), .Y(\reg_file_next[27][8] ) );
  MXI2XL U530 ( .A(n187), .B(n2142), .S0(n2971), .Y(\reg_file_next[27][9] ) );
  MXI2XL U531 ( .A(n188), .B(n2202), .S0(n2971), .Y(\reg_file_next[27][10] )
         );
  MXI2XL U532 ( .A(n189), .B(n2200), .S0(n2971), .Y(\reg_file_next[27][11] )
         );
  MXI2XL U533 ( .A(n190), .B(n2198), .S0(n2971), .Y(\reg_file_next[27][12] )
         );
  MXI2XL U534 ( .A(n191), .B(n2196), .S0(n2971), .Y(\reg_file_next[27][13] )
         );
  MXI2XL U535 ( .A(n192), .B(n2194), .S0(n2971), .Y(\reg_file_next[27][14] )
         );
  MXI2XL U536 ( .A(n193), .B(n2192), .S0(n2971), .Y(\reg_file_next[27][15] )
         );
  MXI2XL U537 ( .A(n194), .B(n2190), .S0(n2971), .Y(\reg_file_next[27][16] )
         );
  MXI2XL U538 ( .A(n195), .B(n2188), .S0(n2971), .Y(\reg_file_next[27][17] )
         );
  MXI2XL U539 ( .A(n196), .B(n2186), .S0(n2971), .Y(\reg_file_next[27][18] )
         );
  MXI2XL U540 ( .A(n197), .B(n2184), .S0(n2971), .Y(\reg_file_next[27][19] )
         );
  MXI2XL U541 ( .A(n198), .B(n2180), .S0(n2971), .Y(\reg_file_next[27][20] )
         );
  MXI2XL U542 ( .A(n199), .B(n2178), .S0(n2971), .Y(\reg_file_next[27][21] )
         );
  MXI2XL U543 ( .A(n200), .B(n2176), .S0(n2971), .Y(\reg_file_next[27][22] )
         );
  MXI2XL U544 ( .A(n201), .B(n2174), .S0(n2971), .Y(\reg_file_next[27][23] )
         );
  MXI2XL U545 ( .A(n202), .B(n2172), .S0(n2971), .Y(\reg_file_next[27][24] )
         );
  MXI2XL U546 ( .A(n203), .B(n2170), .S0(n2971), .Y(\reg_file_next[27][25] )
         );
  MXI2XL U547 ( .A(n204), .B(n2168), .S0(n2971), .Y(\reg_file_next[27][26] )
         );
  MXI2XL U548 ( .A(n205), .B(n2166), .S0(n2971), .Y(\reg_file_next[27][27] )
         );
  MXI2XL U549 ( .A(n206), .B(n2164), .S0(n2971), .Y(\reg_file_next[27][28] )
         );
  MXI2XL U550 ( .A(n207), .B(n2162), .S0(n2971), .Y(\reg_file_next[27][29] )
         );
  MXI2XL U551 ( .A(n208), .B(n2158), .S0(n2971), .Y(\reg_file_next[27][30] )
         );
  MXI2XL U552 ( .A(n209), .B(n2156), .S0(n2971), .Y(\reg_file_next[27][31] )
         );
  MXI2XL U553 ( .A(n1906), .B(n2204), .S0(n2962), .Y(\reg_file_next[6][0] ) );
  MXI2XL U554 ( .A(n2034), .B(n2204), .S0(n2968), .Y(\reg_file_next[2][0] ) );
  MXI2XL U555 ( .A(n1650), .B(n2204), .S0(n2985), .Y(\reg_file_next[14][0] )
         );
  MXI2XL U556 ( .A(n1778), .B(n2204), .S0(n2989), .Y(\reg_file_next[10][0] )
         );
  MXI2XL U557 ( .A(n1394), .B(n2204), .S0(n2976), .Y(\reg_file_next[22][0] )
         );
  MXI2XL U558 ( .A(n1522), .B(n2204), .S0(n2981), .Y(\reg_file_next[18][0] )
         );
  MXI2XL U559 ( .A(n82), .B(n2204), .S0(n2967), .Y(\reg_file_next[30][0] ) );
  MXI2XL U560 ( .A(n1907), .B(n2182), .S0(n2962), .Y(\reg_file_next[6][1] ) );
  MXI2XL U561 ( .A(n2035), .B(n2182), .S0(n2968), .Y(\reg_file_next[2][1] ) );
  MXI2XL U562 ( .A(n1651), .B(n2182), .S0(n2985), .Y(\reg_file_next[14][1] )
         );
  MXI2XL U563 ( .A(n1779), .B(n2182), .S0(n2989), .Y(\reg_file_next[10][1] )
         );
  MXI2XL U564 ( .A(n1395), .B(n2182), .S0(n2976), .Y(\reg_file_next[22][1] )
         );
  MXI2XL U565 ( .A(n1523), .B(n2182), .S0(n2981), .Y(\reg_file_next[18][1] )
         );
  MXI2XL U566 ( .A(n83), .B(n2182), .S0(n2967), .Y(\reg_file_next[30][1] ) );
  MXI2XL U567 ( .A(n1908), .B(n2160), .S0(n2962), .Y(\reg_file_next[6][2] ) );
  MXI2XL U568 ( .A(n2036), .B(n2160), .S0(n2968), .Y(\reg_file_next[2][2] ) );
  MXI2XL U569 ( .A(n1652), .B(n2160), .S0(n2985), .Y(\reg_file_next[14][2] )
         );
  MXI2XL U570 ( .A(n1780), .B(n2160), .S0(n2989), .Y(\reg_file_next[10][2] )
         );
  MXI2XL U571 ( .A(n1396), .B(n2160), .S0(n2976), .Y(\reg_file_next[22][2] )
         );
  MXI2XL U572 ( .A(n1524), .B(n2160), .S0(n2981), .Y(\reg_file_next[18][2] )
         );
  MXI2XL U573 ( .A(n84), .B(n2160), .S0(n2967), .Y(\reg_file_next[30][2] ) );
  MXI2XL U574 ( .A(n1909), .B(n2154), .S0(n2962), .Y(\reg_file_next[6][3] ) );
  MXI2XL U575 ( .A(n2037), .B(n2154), .S0(n2968), .Y(\reg_file_next[2][3] ) );
  MXI2XL U576 ( .A(n1653), .B(n2154), .S0(n2985), .Y(\reg_file_next[14][3] )
         );
  MXI2XL U577 ( .A(n1781), .B(n2154), .S0(n2989), .Y(\reg_file_next[10][3] )
         );
  MXI2XL U578 ( .A(n1397), .B(n2154), .S0(n2976), .Y(\reg_file_next[22][3] )
         );
  MXI2XL U579 ( .A(n1525), .B(n2154), .S0(n2981), .Y(\reg_file_next[18][3] )
         );
  MXI2XL U580 ( .A(n85), .B(n2154), .S0(n2967), .Y(\reg_file_next[30][3] ) );
  MXI2XL U581 ( .A(n1910), .B(n2152), .S0(n2962), .Y(\reg_file_next[6][4] ) );
  MXI2XL U582 ( .A(n2038), .B(n2152), .S0(n2968), .Y(\reg_file_next[2][4] ) );
  MXI2XL U583 ( .A(n1654), .B(n2152), .S0(n2985), .Y(\reg_file_next[14][4] )
         );
  MXI2XL U584 ( .A(n1782), .B(n2152), .S0(n2989), .Y(\reg_file_next[10][4] )
         );
  MXI2XL U585 ( .A(n1398), .B(n2152), .S0(n2976), .Y(\reg_file_next[22][4] )
         );
  MXI2XL U586 ( .A(n1526), .B(n2152), .S0(n2981), .Y(\reg_file_next[18][4] )
         );
  MXI2XL U587 ( .A(n86), .B(n2152), .S0(n2967), .Y(\reg_file_next[30][4] ) );
  MXI2XL U588 ( .A(n1911), .B(n2150), .S0(n2962), .Y(\reg_file_next[6][5] ) );
  MXI2XL U589 ( .A(n2039), .B(n2150), .S0(n2968), .Y(\reg_file_next[2][5] ) );
  MXI2XL U590 ( .A(n1655), .B(n2150), .S0(n2985), .Y(\reg_file_next[14][5] )
         );
  MXI2XL U591 ( .A(n1783), .B(n2150), .S0(n2989), .Y(\reg_file_next[10][5] )
         );
  MXI2XL U592 ( .A(n1399), .B(n2150), .S0(n2976), .Y(\reg_file_next[22][5] )
         );
  MXI2XL U593 ( .A(n1527), .B(n2150), .S0(n2981), .Y(\reg_file_next[18][5] )
         );
  MXI2XL U594 ( .A(n87), .B(n2150), .S0(n2967), .Y(\reg_file_next[30][5] ) );
  MXI2XL U595 ( .A(n1912), .B(n2148), .S0(n2962), .Y(\reg_file_next[6][6] ) );
  MXI2XL U596 ( .A(n2040), .B(n2148), .S0(n2968), .Y(\reg_file_next[2][6] ) );
  MXI2XL U597 ( .A(n1656), .B(n2148), .S0(n2985), .Y(\reg_file_next[14][6] )
         );
  MXI2XL U598 ( .A(n1784), .B(n2148), .S0(n2989), .Y(\reg_file_next[10][6] )
         );
  MXI2XL U599 ( .A(n1400), .B(n2148), .S0(n2976), .Y(\reg_file_next[22][6] )
         );
  MXI2XL U600 ( .A(n1528), .B(n2148), .S0(n2981), .Y(\reg_file_next[18][6] )
         );
  MXI2XL U601 ( .A(n88), .B(n2148), .S0(n2967), .Y(\reg_file_next[30][6] ) );
  MXI2XL U602 ( .A(n1913), .B(n2146), .S0(n2962), .Y(\reg_file_next[6][7] ) );
  MXI2XL U603 ( .A(n2041), .B(n2146), .S0(n2968), .Y(\reg_file_next[2][7] ) );
  MXI2XL U604 ( .A(n1657), .B(n2146), .S0(n2985), .Y(\reg_file_next[14][7] )
         );
  MXI2XL U605 ( .A(n1785), .B(n2146), .S0(n2989), .Y(\reg_file_next[10][7] )
         );
  MXI2XL U606 ( .A(n1401), .B(n2146), .S0(n2976), .Y(\reg_file_next[22][7] )
         );
  MXI2XL U607 ( .A(n1529), .B(n2146), .S0(n2981), .Y(\reg_file_next[18][7] )
         );
  MXI2XL U608 ( .A(n89), .B(n2146), .S0(n2967), .Y(\reg_file_next[30][7] ) );
  MXI2XL U609 ( .A(n1914), .B(n2144), .S0(n2962), .Y(\reg_file_next[6][8] ) );
  MXI2XL U610 ( .A(n2042), .B(n2144), .S0(n2968), .Y(\reg_file_next[2][8] ) );
  MXI2XL U611 ( .A(n1658), .B(n2144), .S0(n2985), .Y(\reg_file_next[14][8] )
         );
  MXI2XL U612 ( .A(n1786), .B(n2144), .S0(n2989), .Y(\reg_file_next[10][8] )
         );
  MXI2XL U613 ( .A(n1402), .B(n2144), .S0(n2976), .Y(\reg_file_next[22][8] )
         );
  MXI2XL U614 ( .A(n1530), .B(n2144), .S0(n2981), .Y(\reg_file_next[18][8] )
         );
  MXI2XL U615 ( .A(n90), .B(n2144), .S0(n2967), .Y(\reg_file_next[30][8] ) );
  MXI2XL U616 ( .A(n1915), .B(n2142), .S0(n2962), .Y(\reg_file_next[6][9] ) );
  MXI2XL U617 ( .A(n2043), .B(n2142), .S0(n2968), .Y(\reg_file_next[2][9] ) );
  MXI2XL U618 ( .A(n1659), .B(n2142), .S0(n2985), .Y(\reg_file_next[14][9] )
         );
  MXI2XL U619 ( .A(n1787), .B(n2142), .S0(n2989), .Y(\reg_file_next[10][9] )
         );
  MXI2XL U620 ( .A(n1403), .B(n2142), .S0(n2976), .Y(\reg_file_next[22][9] )
         );
  MXI2XL U621 ( .A(n1531), .B(n2142), .S0(n2981), .Y(\reg_file_next[18][9] )
         );
  MXI2XL U622 ( .A(n91), .B(n2142), .S0(n2967), .Y(\reg_file_next[30][9] ) );
  MXI2XL U623 ( .A(n1916), .B(n2202), .S0(n2962), .Y(\reg_file_next[6][10] )
         );
  MXI2XL U624 ( .A(n2044), .B(n2202), .S0(n2968), .Y(\reg_file_next[2][10] )
         );
  MXI2XL U625 ( .A(n1660), .B(n2202), .S0(n2985), .Y(\reg_file_next[14][10] )
         );
  MXI2XL U626 ( .A(n1788), .B(n2202), .S0(n2989), .Y(\reg_file_next[10][10] )
         );
  MXI2XL U627 ( .A(n1404), .B(n2202), .S0(n2976), .Y(\reg_file_next[22][10] )
         );
  MXI2XL U628 ( .A(n1532), .B(n2202), .S0(n2981), .Y(\reg_file_next[18][10] )
         );
  MXI2XL U629 ( .A(n92), .B(n2202), .S0(n2967), .Y(\reg_file_next[30][10] ) );
  MXI2XL U630 ( .A(n1917), .B(n2200), .S0(n2962), .Y(\reg_file_next[6][11] )
         );
  MXI2XL U631 ( .A(n2045), .B(n2200), .S0(n2968), .Y(\reg_file_next[2][11] )
         );
  MXI2XL U632 ( .A(n1661), .B(n2200), .S0(n2985), .Y(\reg_file_next[14][11] )
         );
  MXI2XL U633 ( .A(n1789), .B(n2200), .S0(n2989), .Y(\reg_file_next[10][11] )
         );
  MXI2XL U634 ( .A(n1405), .B(n2200), .S0(n2976), .Y(\reg_file_next[22][11] )
         );
  MXI2XL U635 ( .A(n1533), .B(n2200), .S0(n2981), .Y(\reg_file_next[18][11] )
         );
  MXI2XL U636 ( .A(n93), .B(n2200), .S0(n2967), .Y(\reg_file_next[30][11] ) );
  MXI2XL U637 ( .A(n1918), .B(n2198), .S0(n2962), .Y(\reg_file_next[6][12] )
         );
  MXI2XL U638 ( .A(n2046), .B(n2198), .S0(n2968), .Y(\reg_file_next[2][12] )
         );
  MXI2XL U639 ( .A(n1662), .B(n2198), .S0(n2985), .Y(\reg_file_next[14][12] )
         );
  MXI2XL U640 ( .A(n1790), .B(n2198), .S0(n2989), .Y(\reg_file_next[10][12] )
         );
  MXI2XL U641 ( .A(n1406), .B(n2198), .S0(n2976), .Y(\reg_file_next[22][12] )
         );
  MXI2XL U642 ( .A(n1534), .B(n2198), .S0(n2981), .Y(\reg_file_next[18][12] )
         );
  MXI2XL U643 ( .A(n94), .B(n2198), .S0(n2967), .Y(\reg_file_next[30][12] ) );
  MXI2XL U644 ( .A(n1919), .B(n2196), .S0(n2962), .Y(\reg_file_next[6][13] )
         );
  MXI2XL U645 ( .A(n2047), .B(n2196), .S0(n2968), .Y(\reg_file_next[2][13] )
         );
  MXI2XL U646 ( .A(n1663), .B(n2196), .S0(n2985), .Y(\reg_file_next[14][13] )
         );
  MXI2XL U647 ( .A(n1791), .B(n2196), .S0(n2989), .Y(\reg_file_next[10][13] )
         );
  MXI2XL U648 ( .A(n1407), .B(n2196), .S0(n2976), .Y(\reg_file_next[22][13] )
         );
  MXI2XL U649 ( .A(n1535), .B(n2196), .S0(n2981), .Y(\reg_file_next[18][13] )
         );
  MXI2XL U650 ( .A(n95), .B(n2196), .S0(n2967), .Y(\reg_file_next[30][13] ) );
  MXI2XL U651 ( .A(n1920), .B(n2194), .S0(n2962), .Y(\reg_file_next[6][14] )
         );
  MXI2XL U652 ( .A(n2048), .B(n2194), .S0(n2968), .Y(\reg_file_next[2][14] )
         );
  MXI2XL U653 ( .A(n1664), .B(n2194), .S0(n2985), .Y(\reg_file_next[14][14] )
         );
  MXI2XL U654 ( .A(n1792), .B(n2194), .S0(n2989), .Y(\reg_file_next[10][14] )
         );
  MXI2XL U655 ( .A(n1408), .B(n2194), .S0(n2976), .Y(\reg_file_next[22][14] )
         );
  MXI2XL U656 ( .A(n1536), .B(n2194), .S0(n2981), .Y(\reg_file_next[18][14] )
         );
  MXI2XL U657 ( .A(n96), .B(n2194), .S0(n2967), .Y(\reg_file_next[30][14] ) );
  MXI2XL U658 ( .A(n1921), .B(n2192), .S0(n2962), .Y(\reg_file_next[6][15] )
         );
  MXI2XL U659 ( .A(n2049), .B(n2192), .S0(n2968), .Y(\reg_file_next[2][15] )
         );
  MXI2XL U660 ( .A(n1665), .B(n2192), .S0(n2985), .Y(\reg_file_next[14][15] )
         );
  MXI2XL U661 ( .A(n1793), .B(n2192), .S0(n2989), .Y(\reg_file_next[10][15] )
         );
  MXI2XL U662 ( .A(n1409), .B(n2192), .S0(n2976), .Y(\reg_file_next[22][15] )
         );
  MXI2XL U663 ( .A(n1537), .B(n2192), .S0(n2981), .Y(\reg_file_next[18][15] )
         );
  MXI2XL U664 ( .A(n97), .B(n2192), .S0(n2967), .Y(\reg_file_next[30][15] ) );
  MXI2XL U665 ( .A(n1922), .B(n2190), .S0(n2962), .Y(\reg_file_next[6][16] )
         );
  MXI2XL U666 ( .A(n2050), .B(n2190), .S0(n2968), .Y(\reg_file_next[2][16] )
         );
  MXI2XL U667 ( .A(n1666), .B(n2190), .S0(n2985), .Y(\reg_file_next[14][16] )
         );
  MXI2XL U668 ( .A(n1794), .B(n2190), .S0(n2989), .Y(\reg_file_next[10][16] )
         );
  MXI2XL U669 ( .A(n1410), .B(n2190), .S0(n2976), .Y(\reg_file_next[22][16] )
         );
  MXI2XL U670 ( .A(n1538), .B(n2190), .S0(n2981), .Y(\reg_file_next[18][16] )
         );
  MXI2XL U671 ( .A(n98), .B(n2190), .S0(n2967), .Y(\reg_file_next[30][16] ) );
  MXI2XL U672 ( .A(n1923), .B(n2188), .S0(n2962), .Y(\reg_file_next[6][17] )
         );
  MXI2XL U673 ( .A(n2051), .B(n2188), .S0(n2968), .Y(\reg_file_next[2][17] )
         );
  MXI2XL U674 ( .A(n1667), .B(n2188), .S0(n2985), .Y(\reg_file_next[14][17] )
         );
  MXI2XL U675 ( .A(n1795), .B(n2188), .S0(n2989), .Y(\reg_file_next[10][17] )
         );
  MXI2XL U676 ( .A(n1411), .B(n2188), .S0(n2976), .Y(\reg_file_next[22][17] )
         );
  MXI2XL U677 ( .A(n1539), .B(n2188), .S0(n2981), .Y(\reg_file_next[18][17] )
         );
  MXI2XL U678 ( .A(n99), .B(n2188), .S0(n2967), .Y(\reg_file_next[30][17] ) );
  MXI2XL U679 ( .A(n1924), .B(n2186), .S0(n2962), .Y(\reg_file_next[6][18] )
         );
  MXI2XL U680 ( .A(n2052), .B(n2186), .S0(n2968), .Y(\reg_file_next[2][18] )
         );
  MXI2XL U681 ( .A(n1668), .B(n2186), .S0(n2985), .Y(\reg_file_next[14][18] )
         );
  MXI2XL U682 ( .A(n1796), .B(n2186), .S0(n2989), .Y(\reg_file_next[10][18] )
         );
  MXI2XL U683 ( .A(n1412), .B(n2186), .S0(n2976), .Y(\reg_file_next[22][18] )
         );
  MXI2XL U684 ( .A(n1540), .B(n2186), .S0(n2981), .Y(\reg_file_next[18][18] )
         );
  MXI2XL U685 ( .A(n100), .B(n2186), .S0(n2967), .Y(\reg_file_next[30][18] )
         );
  MXI2XL U686 ( .A(n1925), .B(n2184), .S0(n2962), .Y(\reg_file_next[6][19] )
         );
  MXI2XL U687 ( .A(n2053), .B(n2184), .S0(n2968), .Y(\reg_file_next[2][19] )
         );
  MXI2XL U688 ( .A(n1669), .B(n2184), .S0(n2985), .Y(\reg_file_next[14][19] )
         );
  MXI2XL U689 ( .A(n1797), .B(n2184), .S0(n2989), .Y(\reg_file_next[10][19] )
         );
  MXI2XL U690 ( .A(n1413), .B(n2184), .S0(n2976), .Y(\reg_file_next[22][19] )
         );
  MXI2XL U691 ( .A(n1541), .B(n2184), .S0(n2981), .Y(\reg_file_next[18][19] )
         );
  MXI2XL U692 ( .A(n101), .B(n2184), .S0(n2967), .Y(\reg_file_next[30][19] )
         );
  MXI2XL U693 ( .A(n1926), .B(n2180), .S0(n2962), .Y(\reg_file_next[6][20] )
         );
  MXI2XL U694 ( .A(n2054), .B(n2180), .S0(n2968), .Y(\reg_file_next[2][20] )
         );
  MXI2XL U695 ( .A(n1670), .B(n2180), .S0(n2985), .Y(\reg_file_next[14][20] )
         );
  MXI2XL U696 ( .A(n1798), .B(n2180), .S0(n2989), .Y(\reg_file_next[10][20] )
         );
  MXI2XL U697 ( .A(n1414), .B(n2180), .S0(n2976), .Y(\reg_file_next[22][20] )
         );
  MXI2XL U698 ( .A(n1542), .B(n2180), .S0(n2981), .Y(\reg_file_next[18][20] )
         );
  MXI2XL U699 ( .A(n102), .B(n2180), .S0(n2967), .Y(\reg_file_next[30][20] )
         );
  MXI2XL U700 ( .A(n1927), .B(n2178), .S0(n2962), .Y(\reg_file_next[6][21] )
         );
  MXI2XL U701 ( .A(n2055), .B(n2178), .S0(n2968), .Y(\reg_file_next[2][21] )
         );
  MXI2XL U702 ( .A(n1671), .B(n2178), .S0(n2985), .Y(\reg_file_next[14][21] )
         );
  MXI2XL U703 ( .A(n1799), .B(n2178), .S0(n2989), .Y(\reg_file_next[10][21] )
         );
  MXI2XL U704 ( .A(n1415), .B(n2178), .S0(n2976), .Y(\reg_file_next[22][21] )
         );
  MXI2XL U705 ( .A(n1543), .B(n2178), .S0(n2981), .Y(\reg_file_next[18][21] )
         );
  MXI2XL U706 ( .A(n103), .B(n2178), .S0(n2967), .Y(\reg_file_next[30][21] )
         );
  MXI2XL U707 ( .A(n1928), .B(n2176), .S0(n2962), .Y(\reg_file_next[6][22] )
         );
  MXI2XL U708 ( .A(n2056), .B(n2176), .S0(n2968), .Y(\reg_file_next[2][22] )
         );
  MXI2XL U709 ( .A(n1672), .B(n2176), .S0(n2985), .Y(\reg_file_next[14][22] )
         );
  MXI2XL U710 ( .A(n1800), .B(n2176), .S0(n2989), .Y(\reg_file_next[10][22] )
         );
  MXI2XL U711 ( .A(n1416), .B(n2176), .S0(n2976), .Y(\reg_file_next[22][22] )
         );
  MXI2XL U712 ( .A(n1544), .B(n2176), .S0(n2981), .Y(\reg_file_next[18][22] )
         );
  MXI2XL U713 ( .A(n104), .B(n2176), .S0(n2967), .Y(\reg_file_next[30][22] )
         );
  MXI2XL U714 ( .A(n1929), .B(n2174), .S0(n2962), .Y(\reg_file_next[6][23] )
         );
  MXI2XL U715 ( .A(n2057), .B(n2174), .S0(n2968), .Y(\reg_file_next[2][23] )
         );
  MXI2XL U716 ( .A(n1673), .B(n2174), .S0(n2985), .Y(\reg_file_next[14][23] )
         );
  MXI2XL U717 ( .A(n1801), .B(n2174), .S0(n2989), .Y(\reg_file_next[10][23] )
         );
  MXI2XL U718 ( .A(n1417), .B(n2174), .S0(n2976), .Y(\reg_file_next[22][23] )
         );
  MXI2XL U719 ( .A(n1545), .B(n2174), .S0(n2981), .Y(\reg_file_next[18][23] )
         );
  MXI2XL U720 ( .A(n105), .B(n2174), .S0(n2967), .Y(\reg_file_next[30][23] )
         );
  MXI2XL U721 ( .A(n1930), .B(n2172), .S0(n2962), .Y(\reg_file_next[6][24] )
         );
  MXI2XL U722 ( .A(n2058), .B(n2172), .S0(n2968), .Y(\reg_file_next[2][24] )
         );
  MXI2XL U723 ( .A(n1674), .B(n2172), .S0(n2985), .Y(\reg_file_next[14][24] )
         );
  MXI2XL U724 ( .A(n1802), .B(n2172), .S0(n2989), .Y(\reg_file_next[10][24] )
         );
  MXI2XL U725 ( .A(n1418), .B(n2172), .S0(n2976), .Y(\reg_file_next[22][24] )
         );
  MXI2XL U726 ( .A(n1546), .B(n2172), .S0(n2981), .Y(\reg_file_next[18][24] )
         );
  MXI2XL U727 ( .A(n106), .B(n2172), .S0(n2967), .Y(\reg_file_next[30][24] )
         );
  MXI2XL U728 ( .A(n1931), .B(n2170), .S0(n2962), .Y(\reg_file_next[6][25] )
         );
  MXI2XL U729 ( .A(n2059), .B(n2170), .S0(n2968), .Y(\reg_file_next[2][25] )
         );
  MXI2XL U730 ( .A(n1675), .B(n2170), .S0(n2985), .Y(\reg_file_next[14][25] )
         );
  MXI2XL U731 ( .A(n1803), .B(n2170), .S0(n2989), .Y(\reg_file_next[10][25] )
         );
  MXI2XL U732 ( .A(n1419), .B(n2170), .S0(n2976), .Y(\reg_file_next[22][25] )
         );
  MXI2XL U733 ( .A(n1547), .B(n2170), .S0(n2981), .Y(\reg_file_next[18][25] )
         );
  MXI2XL U734 ( .A(n107), .B(n2170), .S0(n2967), .Y(\reg_file_next[30][25] )
         );
  MXI2XL U735 ( .A(n1932), .B(n2168), .S0(n2962), .Y(\reg_file_next[6][26] )
         );
  MXI2XL U736 ( .A(n2060), .B(n2168), .S0(n2968), .Y(\reg_file_next[2][26] )
         );
  MXI2XL U737 ( .A(n1676), .B(n2168), .S0(n2985), .Y(\reg_file_next[14][26] )
         );
  MXI2XL U738 ( .A(n1804), .B(n2168), .S0(n2989), .Y(\reg_file_next[10][26] )
         );
  MXI2XL U739 ( .A(n1420), .B(n2168), .S0(n2976), .Y(\reg_file_next[22][26] )
         );
  MXI2XL U740 ( .A(n1548), .B(n2168), .S0(n2981), .Y(\reg_file_next[18][26] )
         );
  MXI2XL U741 ( .A(n108), .B(n2168), .S0(n2967), .Y(\reg_file_next[30][26] )
         );
  MXI2XL U742 ( .A(n1933), .B(n2166), .S0(n2962), .Y(\reg_file_next[6][27] )
         );
  MXI2XL U743 ( .A(n2061), .B(n2166), .S0(n2968), .Y(\reg_file_next[2][27] )
         );
  MXI2XL U744 ( .A(n1677), .B(n2166), .S0(n2985), .Y(\reg_file_next[14][27] )
         );
  MXI2XL U745 ( .A(n1805), .B(n2166), .S0(n2989), .Y(\reg_file_next[10][27] )
         );
  MXI2XL U746 ( .A(n1421), .B(n2166), .S0(n2976), .Y(\reg_file_next[22][27] )
         );
  MXI2XL U747 ( .A(n1549), .B(n2166), .S0(n2981), .Y(\reg_file_next[18][27] )
         );
  MXI2XL U748 ( .A(n109), .B(n2166), .S0(n2967), .Y(\reg_file_next[30][27] )
         );
  MXI2XL U749 ( .A(n1934), .B(n2164), .S0(n2962), .Y(\reg_file_next[6][28] )
         );
  MXI2XL U750 ( .A(n2062), .B(n2164), .S0(n2968), .Y(\reg_file_next[2][28] )
         );
  MXI2XL U751 ( .A(n1678), .B(n2164), .S0(n2985), .Y(\reg_file_next[14][28] )
         );
  MXI2XL U752 ( .A(n1806), .B(n2164), .S0(n2989), .Y(\reg_file_next[10][28] )
         );
  MXI2XL U753 ( .A(n1422), .B(n2164), .S0(n2976), .Y(\reg_file_next[22][28] )
         );
  MXI2XL U754 ( .A(n1550), .B(n2164), .S0(n2981), .Y(\reg_file_next[18][28] )
         );
  MXI2XL U755 ( .A(n110), .B(n2164), .S0(n2967), .Y(\reg_file_next[30][28] )
         );
  MXI2XL U756 ( .A(n1935), .B(n2162), .S0(n2962), .Y(\reg_file_next[6][29] )
         );
  MXI2XL U757 ( .A(n2063), .B(n2162), .S0(n2968), .Y(\reg_file_next[2][29] )
         );
  MXI2XL U758 ( .A(n1679), .B(n2162), .S0(n2985), .Y(\reg_file_next[14][29] )
         );
  MXI2XL U759 ( .A(n1807), .B(n2162), .S0(n2989), .Y(\reg_file_next[10][29] )
         );
  MXI2XL U760 ( .A(n1423), .B(n2162), .S0(n2976), .Y(\reg_file_next[22][29] )
         );
  MXI2XL U761 ( .A(n1551), .B(n2162), .S0(n2981), .Y(\reg_file_next[18][29] )
         );
  MXI2XL U762 ( .A(n111), .B(n2162), .S0(n2967), .Y(\reg_file_next[30][29] )
         );
  MXI2XL U763 ( .A(n1936), .B(n2158), .S0(n2962), .Y(\reg_file_next[6][30] )
         );
  MXI2XL U764 ( .A(n2064), .B(n2158), .S0(n2968), .Y(\reg_file_next[2][30] )
         );
  MXI2XL U765 ( .A(n1680), .B(n2158), .S0(n2985), .Y(\reg_file_next[14][30] )
         );
  MXI2XL U766 ( .A(n1808), .B(n2158), .S0(n2989), .Y(\reg_file_next[10][30] )
         );
  MXI2XL U767 ( .A(n1424), .B(n2158), .S0(n2976), .Y(\reg_file_next[22][30] )
         );
  MXI2XL U768 ( .A(n1552), .B(n2158), .S0(n2981), .Y(\reg_file_next[18][30] )
         );
  MXI2XL U769 ( .A(n112), .B(n2158), .S0(n2967), .Y(\reg_file_next[30][30] )
         );
  MXI2XL U770 ( .A(n1937), .B(n2156), .S0(n2962), .Y(\reg_file_next[6][31] )
         );
  MXI2XL U771 ( .A(n2065), .B(n2156), .S0(n2968), .Y(\reg_file_next[2][31] )
         );
  MXI2XL U772 ( .A(n1681), .B(n2156), .S0(n2985), .Y(\reg_file_next[14][31] )
         );
  MXI2XL U773 ( .A(n1809), .B(n2156), .S0(n2989), .Y(\reg_file_next[10][31] )
         );
  MXI2XL U774 ( .A(n1425), .B(n2156), .S0(n2976), .Y(\reg_file_next[22][31] )
         );
  MXI2XL U775 ( .A(n1553), .B(n2156), .S0(n2981), .Y(\reg_file_next[18][31] )
         );
  MXI2XL U776 ( .A(n113), .B(n2156), .S0(n2967), .Y(\reg_file_next[30][31] )
         );
  MXI2XL U777 ( .A(n210), .B(n2204), .S0(n2972), .Y(\reg_file_next[26][0] ) );
  MXI2XL U778 ( .A(n211), .B(n2182), .S0(n2972), .Y(\reg_file_next[26][1] ) );
  MXI2XL U779 ( .A(n212), .B(n2160), .S0(n2972), .Y(\reg_file_next[26][2] ) );
  MXI2XL U780 ( .A(n213), .B(n2154), .S0(n2972), .Y(\reg_file_next[26][3] ) );
  MXI2XL U781 ( .A(n214), .B(n2152), .S0(n2972), .Y(\reg_file_next[26][4] ) );
  MXI2XL U782 ( .A(n215), .B(n2150), .S0(n2972), .Y(\reg_file_next[26][5] ) );
  MXI2XL U783 ( .A(n216), .B(n2148), .S0(n2972), .Y(\reg_file_next[26][6] ) );
  MXI2XL U784 ( .A(n217), .B(n2146), .S0(n2972), .Y(\reg_file_next[26][7] ) );
  MXI2XL U785 ( .A(n218), .B(n2144), .S0(n2972), .Y(\reg_file_next[26][8] ) );
  MXI2XL U786 ( .A(n219), .B(n2142), .S0(n2972), .Y(\reg_file_next[26][9] ) );
  MXI2XL U787 ( .A(n220), .B(n2202), .S0(n2972), .Y(\reg_file_next[26][10] )
         );
  MXI2XL U788 ( .A(n221), .B(n2200), .S0(n2972), .Y(\reg_file_next[26][11] )
         );
  MXI2XL U789 ( .A(n222), .B(n2198), .S0(n2972), .Y(\reg_file_next[26][12] )
         );
  MXI2XL U790 ( .A(n223), .B(n2196), .S0(n2972), .Y(\reg_file_next[26][13] )
         );
  MXI2XL U791 ( .A(n224), .B(n2194), .S0(n2972), .Y(\reg_file_next[26][14] )
         );
  MXI2XL U792 ( .A(n225), .B(n2192), .S0(n2972), .Y(\reg_file_next[26][15] )
         );
  MXI2XL U793 ( .A(n226), .B(n2190), .S0(n2972), .Y(\reg_file_next[26][16] )
         );
  MXI2XL U794 ( .A(n227), .B(n2188), .S0(n2972), .Y(\reg_file_next[26][17] )
         );
  MXI2XL U795 ( .A(n228), .B(n2186), .S0(n2972), .Y(\reg_file_next[26][18] )
         );
  MXI2XL U796 ( .A(n229), .B(n2184), .S0(n2972), .Y(\reg_file_next[26][19] )
         );
  MXI2XL U797 ( .A(n230), .B(n2180), .S0(n2972), .Y(\reg_file_next[26][20] )
         );
  MXI2XL U798 ( .A(n231), .B(n2178), .S0(n2972), .Y(\reg_file_next[26][21] )
         );
  MXI2XL U799 ( .A(n232), .B(n2176), .S0(n2972), .Y(\reg_file_next[26][22] )
         );
  MXI2XL U800 ( .A(n233), .B(n2174), .S0(n2972), .Y(\reg_file_next[26][23] )
         );
  MXI2XL U801 ( .A(n234), .B(n2172), .S0(n2972), .Y(\reg_file_next[26][24] )
         );
  MXI2XL U802 ( .A(n235), .B(n2170), .S0(n2972), .Y(\reg_file_next[26][25] )
         );
  MXI2XL U803 ( .A(n236), .B(n2168), .S0(n2972), .Y(\reg_file_next[26][26] )
         );
  MXI2XL U804 ( .A(n237), .B(n2166), .S0(n2972), .Y(\reg_file_next[26][27] )
         );
  MXI2XL U805 ( .A(n238), .B(n2164), .S0(n2972), .Y(\reg_file_next[26][28] )
         );
  MXI2XL U806 ( .A(n239), .B(n2162), .S0(n2972), .Y(\reg_file_next[26][29] )
         );
  MXI2XL U807 ( .A(n240), .B(n2158), .S0(n2972), .Y(\reg_file_next[26][30] )
         );
  MXI2XL U808 ( .A(n241), .B(n2156), .S0(n2972), .Y(\reg_file_next[26][31] )
         );
  MXI2XL U809 ( .A(n1970), .B(n2204), .S0(n2964), .Y(\reg_file_next[4][0] ) );
  MXI2XL U810 ( .A(n2098), .B(n2204), .S0(n2990), .Y(\reg_file_next[0][0] ) );
  MXI2XL U811 ( .A(n1714), .B(n2204), .S0(n2987), .Y(\reg_file_next[12][0] )
         );
  MXI2XL U812 ( .A(n1842), .B(n2204), .S0(n2960), .Y(\reg_file_next[8][0] ) );
  MXI2XL U813 ( .A(n1458), .B(n2204), .S0(n2978), .Y(\reg_file_next[20][0] )
         );
  MXI2XL U814 ( .A(n1586), .B(n2204), .S0(n2983), .Y(\reg_file_next[16][0] )
         );
  MXI2XL U815 ( .A(n146), .B(n2204), .S0(n2970), .Y(\reg_file_next[28][0] ) );
  MXI2XL U816 ( .A(n1971), .B(n2182), .S0(n2964), .Y(\reg_file_next[4][1] ) );
  MXI2XL U817 ( .A(n2099), .B(n2182), .S0(n2990), .Y(\reg_file_next[0][1] ) );
  MXI2XL U818 ( .A(n1715), .B(n2182), .S0(n2987), .Y(\reg_file_next[12][1] )
         );
  MXI2XL U819 ( .A(n1843), .B(n2182), .S0(n2960), .Y(\reg_file_next[8][1] ) );
  MXI2XL U820 ( .A(n1459), .B(n2182), .S0(n2978), .Y(\reg_file_next[20][1] )
         );
  MXI2XL U821 ( .A(n1587), .B(n2182), .S0(n2983), .Y(\reg_file_next[16][1] )
         );
  MXI2XL U822 ( .A(n147), .B(n2182), .S0(n2970), .Y(\reg_file_next[28][1] ) );
  MXI2XL U823 ( .A(n1972), .B(n2160), .S0(n2964), .Y(\reg_file_next[4][2] ) );
  MXI2XL U824 ( .A(n2100), .B(n2160), .S0(n2990), .Y(\reg_file_next[0][2] ) );
  MXI2XL U825 ( .A(n1716), .B(n2160), .S0(n2987), .Y(\reg_file_next[12][2] )
         );
  MXI2XL U826 ( .A(n1844), .B(n2160), .S0(n2960), .Y(\reg_file_next[8][2] ) );
  MXI2XL U827 ( .A(n1460), .B(n2160), .S0(n2978), .Y(\reg_file_next[20][2] )
         );
  MXI2XL U828 ( .A(n1588), .B(n2160), .S0(n2983), .Y(\reg_file_next[16][2] )
         );
  MXI2XL U829 ( .A(n148), .B(n2160), .S0(n2970), .Y(\reg_file_next[28][2] ) );
  MXI2XL U830 ( .A(n1973), .B(n2154), .S0(n2964), .Y(\reg_file_next[4][3] ) );
  MXI2XL U831 ( .A(n2101), .B(n2154), .S0(n2990), .Y(\reg_file_next[0][3] ) );
  MXI2XL U832 ( .A(n1717), .B(n2154), .S0(n2987), .Y(\reg_file_next[12][3] )
         );
  MXI2XL U833 ( .A(n1845), .B(n2154), .S0(n2960), .Y(\reg_file_next[8][3] ) );
  MXI2XL U834 ( .A(n1461), .B(n2154), .S0(n2978), .Y(\reg_file_next[20][3] )
         );
  MXI2XL U835 ( .A(n1589), .B(n2154), .S0(n2983), .Y(\reg_file_next[16][3] )
         );
  MXI2XL U836 ( .A(n149), .B(n2154), .S0(n2970), .Y(\reg_file_next[28][3] ) );
  MXI2XL U837 ( .A(n1974), .B(n2152), .S0(n2964), .Y(\reg_file_next[4][4] ) );
  MXI2XL U838 ( .A(n2102), .B(n2152), .S0(n2990), .Y(\reg_file_next[0][4] ) );
  MXI2XL U839 ( .A(n1718), .B(n2152), .S0(n2987), .Y(\reg_file_next[12][4] )
         );
  MXI2XL U840 ( .A(n1846), .B(n2152), .S0(n2960), .Y(\reg_file_next[8][4] ) );
  MXI2XL U841 ( .A(n1462), .B(n2152), .S0(n2978), .Y(\reg_file_next[20][4] )
         );
  MXI2XL U842 ( .A(n1590), .B(n2152), .S0(n2983), .Y(\reg_file_next[16][4] )
         );
  MXI2XL U843 ( .A(n150), .B(n2152), .S0(n2970), .Y(\reg_file_next[28][4] ) );
  MXI2XL U844 ( .A(n1975), .B(n2150), .S0(n2964), .Y(\reg_file_next[4][5] ) );
  MXI2XL U845 ( .A(n2103), .B(n2150), .S0(n2990), .Y(\reg_file_next[0][5] ) );
  MXI2XL U846 ( .A(n1719), .B(n2150), .S0(n2987), .Y(\reg_file_next[12][5] )
         );
  MXI2XL U847 ( .A(n1847), .B(n2150), .S0(n2960), .Y(\reg_file_next[8][5] ) );
  MXI2XL U848 ( .A(n1463), .B(n2150), .S0(n2978), .Y(\reg_file_next[20][5] )
         );
  MXI2XL U849 ( .A(n1591), .B(n2150), .S0(n2983), .Y(\reg_file_next[16][5] )
         );
  MXI2XL U850 ( .A(n151), .B(n2150), .S0(n2970), .Y(\reg_file_next[28][5] ) );
  MXI2XL U851 ( .A(n1976), .B(n2148), .S0(n2964), .Y(\reg_file_next[4][6] ) );
  MXI2XL U852 ( .A(n2104), .B(n2148), .S0(n2990), .Y(\reg_file_next[0][6] ) );
  MXI2XL U853 ( .A(n1720), .B(n2148), .S0(n2987), .Y(\reg_file_next[12][6] )
         );
  MXI2XL U854 ( .A(n1848), .B(n2148), .S0(n2960), .Y(\reg_file_next[8][6] ) );
  MXI2XL U855 ( .A(n1464), .B(n2148), .S0(n2978), .Y(\reg_file_next[20][6] )
         );
  MXI2XL U856 ( .A(n1592), .B(n2148), .S0(n2983), .Y(\reg_file_next[16][6] )
         );
  MXI2XL U857 ( .A(n152), .B(n2148), .S0(n2970), .Y(\reg_file_next[28][6] ) );
  MXI2XL U858 ( .A(n1977), .B(n2146), .S0(n2964), .Y(\reg_file_next[4][7] ) );
  MXI2XL U859 ( .A(n2105), .B(n2146), .S0(n2990), .Y(\reg_file_next[0][7] ) );
  MXI2XL U860 ( .A(n1721), .B(n2146), .S0(n2987), .Y(\reg_file_next[12][7] )
         );
  MXI2XL U861 ( .A(n1849), .B(n2146), .S0(n2960), .Y(\reg_file_next[8][7] ) );
  MXI2XL U862 ( .A(n1465), .B(n2146), .S0(n2978), .Y(\reg_file_next[20][7] )
         );
  MXI2XL U863 ( .A(n1593), .B(n2146), .S0(n2983), .Y(\reg_file_next[16][7] )
         );
  MXI2XL U864 ( .A(n153), .B(n2146), .S0(n2970), .Y(\reg_file_next[28][7] ) );
  MXI2XL U865 ( .A(n1978), .B(n2144), .S0(n2964), .Y(\reg_file_next[4][8] ) );
  MXI2XL U866 ( .A(n2106), .B(n2144), .S0(n2990), .Y(\reg_file_next[0][8] ) );
  MXI2XL U867 ( .A(n1722), .B(n2144), .S0(n2987), .Y(\reg_file_next[12][8] )
         );
  MXI2XL U868 ( .A(n1850), .B(n2144), .S0(n2960), .Y(\reg_file_next[8][8] ) );
  MXI2XL U869 ( .A(n1466), .B(n2144), .S0(n2978), .Y(\reg_file_next[20][8] )
         );
  MXI2XL U870 ( .A(n1594), .B(n2144), .S0(n2983), .Y(\reg_file_next[16][8] )
         );
  MXI2XL U871 ( .A(n154), .B(n2144), .S0(n2970), .Y(\reg_file_next[28][8] ) );
  MXI2XL U872 ( .A(n1979), .B(n2142), .S0(n2964), .Y(\reg_file_next[4][9] ) );
  MXI2XL U873 ( .A(n2107), .B(n2142), .S0(n2990), .Y(\reg_file_next[0][9] ) );
  MXI2XL U874 ( .A(n1723), .B(n2142), .S0(n2987), .Y(\reg_file_next[12][9] )
         );
  MXI2XL U875 ( .A(n1851), .B(n2142), .S0(n2960), .Y(\reg_file_next[8][9] ) );
  MXI2XL U876 ( .A(n1467), .B(n2142), .S0(n2978), .Y(\reg_file_next[20][9] )
         );
  MXI2XL U877 ( .A(n1595), .B(n2142), .S0(n2983), .Y(\reg_file_next[16][9] )
         );
  MXI2XL U878 ( .A(n155), .B(n2142), .S0(n2970), .Y(\reg_file_next[28][9] ) );
  MXI2XL U879 ( .A(n1980), .B(n2202), .S0(n2964), .Y(\reg_file_next[4][10] )
         );
  MXI2XL U880 ( .A(n2108), .B(n2202), .S0(n2990), .Y(\reg_file_next[0][10] )
         );
  MXI2XL U881 ( .A(n1724), .B(n2202), .S0(n2987), .Y(\reg_file_next[12][10] )
         );
  MXI2XL U882 ( .A(n1852), .B(n2202), .S0(n2960), .Y(\reg_file_next[8][10] )
         );
  MXI2XL U883 ( .A(n1468), .B(n2202), .S0(n2978), .Y(\reg_file_next[20][10] )
         );
  MXI2XL U884 ( .A(n1596), .B(n2202), .S0(n2983), .Y(\reg_file_next[16][10] )
         );
  MXI2XL U885 ( .A(n156), .B(n2202), .S0(n2970), .Y(\reg_file_next[28][10] )
         );
  MXI2XL U886 ( .A(n1981), .B(n2200), .S0(n2964), .Y(\reg_file_next[4][11] )
         );
  MXI2XL U887 ( .A(n2109), .B(n2200), .S0(n2990), .Y(\reg_file_next[0][11] )
         );
  MXI2XL U888 ( .A(n1725), .B(n2200), .S0(n2987), .Y(\reg_file_next[12][11] )
         );
  MXI2XL U889 ( .A(n1853), .B(n2200), .S0(n2960), .Y(\reg_file_next[8][11] )
         );
  MXI2XL U890 ( .A(n1469), .B(n2200), .S0(n2978), .Y(\reg_file_next[20][11] )
         );
  MXI2XL U891 ( .A(n1597), .B(n2200), .S0(n2983), .Y(\reg_file_next[16][11] )
         );
  MXI2XL U892 ( .A(n157), .B(n2200), .S0(n2970), .Y(\reg_file_next[28][11] )
         );
  MXI2XL U893 ( .A(n1982), .B(n2198), .S0(n2964), .Y(\reg_file_next[4][12] )
         );
  MXI2XL U894 ( .A(n2110), .B(n2198), .S0(n2990), .Y(\reg_file_next[0][12] )
         );
  MXI2XL U895 ( .A(n1726), .B(n2198), .S0(n2987), .Y(\reg_file_next[12][12] )
         );
  MXI2XL U896 ( .A(n1854), .B(n2198), .S0(n2960), .Y(\reg_file_next[8][12] )
         );
  MXI2XL U897 ( .A(n1470), .B(n2198), .S0(n2978), .Y(\reg_file_next[20][12] )
         );
  MXI2XL U898 ( .A(n1598), .B(n2198), .S0(n2983), .Y(\reg_file_next[16][12] )
         );
  MXI2XL U899 ( .A(n158), .B(n2198), .S0(n2970), .Y(\reg_file_next[28][12] )
         );
  MXI2XL U900 ( .A(n1983), .B(n2196), .S0(n2964), .Y(\reg_file_next[4][13] )
         );
  MXI2XL U901 ( .A(n2111), .B(n2196), .S0(n2990), .Y(\reg_file_next[0][13] )
         );
  MXI2XL U902 ( .A(n1727), .B(n2196), .S0(n2987), .Y(\reg_file_next[12][13] )
         );
  MXI2XL U903 ( .A(n1855), .B(n2196), .S0(n2960), .Y(\reg_file_next[8][13] )
         );
  MXI2XL U904 ( .A(n1471), .B(n2196), .S0(n2978), .Y(\reg_file_next[20][13] )
         );
  MXI2XL U905 ( .A(n1599), .B(n2196), .S0(n2983), .Y(\reg_file_next[16][13] )
         );
  MXI2XL U906 ( .A(n159), .B(n2196), .S0(n2970), .Y(\reg_file_next[28][13] )
         );
  MXI2XL U907 ( .A(n1984), .B(n2194), .S0(n2964), .Y(\reg_file_next[4][14] )
         );
  MXI2XL U908 ( .A(n2112), .B(n2194), .S0(n2990), .Y(\reg_file_next[0][14] )
         );
  MXI2XL U909 ( .A(n1728), .B(n2194), .S0(n2987), .Y(\reg_file_next[12][14] )
         );
  MXI2XL U910 ( .A(n1856), .B(n2194), .S0(n2960), .Y(\reg_file_next[8][14] )
         );
  MXI2XL U911 ( .A(n1472), .B(n2194), .S0(n2978), .Y(\reg_file_next[20][14] )
         );
  MXI2XL U912 ( .A(n1600), .B(n2194), .S0(n2983), .Y(\reg_file_next[16][14] )
         );
  MXI2XL U913 ( .A(n160), .B(n2194), .S0(n2970), .Y(\reg_file_next[28][14] )
         );
  MXI2XL U914 ( .A(n1985), .B(n2192), .S0(n2964), .Y(\reg_file_next[4][15] )
         );
  MXI2XL U915 ( .A(n2113), .B(n2192), .S0(n2990), .Y(\reg_file_next[0][15] )
         );
  MXI2XL U916 ( .A(n1729), .B(n2192), .S0(n2987), .Y(\reg_file_next[12][15] )
         );
  MXI2XL U917 ( .A(n1857), .B(n2192), .S0(n2960), .Y(\reg_file_next[8][15] )
         );
  MXI2XL U918 ( .A(n1473), .B(n2192), .S0(n2978), .Y(\reg_file_next[20][15] )
         );
  MXI2XL U919 ( .A(n1601), .B(n2192), .S0(n2983), .Y(\reg_file_next[16][15] )
         );
  MXI2XL U920 ( .A(n161), .B(n2192), .S0(n2970), .Y(\reg_file_next[28][15] )
         );
  MXI2XL U921 ( .A(n1986), .B(n2190), .S0(n2964), .Y(\reg_file_next[4][16] )
         );
  MXI2XL U922 ( .A(n2114), .B(n2190), .S0(n2990), .Y(\reg_file_next[0][16] )
         );
  MXI2XL U923 ( .A(n1730), .B(n2190), .S0(n2987), .Y(\reg_file_next[12][16] )
         );
  MXI2XL U924 ( .A(n1858), .B(n2190), .S0(n2960), .Y(\reg_file_next[8][16] )
         );
  MXI2XL U925 ( .A(n1474), .B(n2190), .S0(n2978), .Y(\reg_file_next[20][16] )
         );
  MXI2XL U926 ( .A(n1602), .B(n2190), .S0(n2983), .Y(\reg_file_next[16][16] )
         );
  MXI2XL U927 ( .A(n162), .B(n2190), .S0(n2970), .Y(\reg_file_next[28][16] )
         );
  MXI2XL U928 ( .A(n1987), .B(n2188), .S0(n2964), .Y(\reg_file_next[4][17] )
         );
  MXI2XL U929 ( .A(n2115), .B(n2188), .S0(n2990), .Y(\reg_file_next[0][17] )
         );
  MXI2XL U930 ( .A(n1731), .B(n2188), .S0(n2987), .Y(\reg_file_next[12][17] )
         );
  MXI2XL U931 ( .A(n1859), .B(n2188), .S0(n2960), .Y(\reg_file_next[8][17] )
         );
  MXI2XL U932 ( .A(n1475), .B(n2188), .S0(n2978), .Y(\reg_file_next[20][17] )
         );
  MXI2XL U933 ( .A(n1603), .B(n2188), .S0(n2983), .Y(\reg_file_next[16][17] )
         );
  MXI2XL U934 ( .A(n163), .B(n2188), .S0(n2970), .Y(\reg_file_next[28][17] )
         );
  MXI2XL U935 ( .A(n1988), .B(n2186), .S0(n2964), .Y(\reg_file_next[4][18] )
         );
  MXI2XL U936 ( .A(n2116), .B(n2186), .S0(n2990), .Y(\reg_file_next[0][18] )
         );
  MXI2XL U937 ( .A(n1732), .B(n2186), .S0(n2987), .Y(\reg_file_next[12][18] )
         );
  MXI2XL U938 ( .A(n1860), .B(n2186), .S0(n2960), .Y(\reg_file_next[8][18] )
         );
  MXI2XL U939 ( .A(n1476), .B(n2186), .S0(n2978), .Y(\reg_file_next[20][18] )
         );
  MXI2XL U940 ( .A(n1604), .B(n2186), .S0(n2983), .Y(\reg_file_next[16][18] )
         );
  MXI2XL U941 ( .A(n164), .B(n2186), .S0(n2970), .Y(\reg_file_next[28][18] )
         );
  MXI2XL U942 ( .A(n1989), .B(n2184), .S0(n2964), .Y(\reg_file_next[4][19] )
         );
  MXI2XL U943 ( .A(n2117), .B(n2184), .S0(n2990), .Y(\reg_file_next[0][19] )
         );
  MXI2XL U944 ( .A(n1733), .B(n2184), .S0(n2987), .Y(\reg_file_next[12][19] )
         );
  MXI2XL U945 ( .A(n1861), .B(n2184), .S0(n2960), .Y(\reg_file_next[8][19] )
         );
  MXI2XL U946 ( .A(n1477), .B(n2184), .S0(n2978), .Y(\reg_file_next[20][19] )
         );
  MXI2XL U947 ( .A(n1605), .B(n2184), .S0(n2983), .Y(\reg_file_next[16][19] )
         );
  MXI2XL U948 ( .A(n165), .B(n2184), .S0(n2970), .Y(\reg_file_next[28][19] )
         );
  MXI2XL U949 ( .A(n1990), .B(n2180), .S0(n2964), .Y(\reg_file_next[4][20] )
         );
  MXI2XL U950 ( .A(n2118), .B(n2180), .S0(n2990), .Y(\reg_file_next[0][20] )
         );
  MXI2XL U951 ( .A(n1734), .B(n2180), .S0(n2987), .Y(\reg_file_next[12][20] )
         );
  MXI2XL U952 ( .A(n1862), .B(n2180), .S0(n2960), .Y(\reg_file_next[8][20] )
         );
  MXI2XL U953 ( .A(n1478), .B(n2180), .S0(n2978), .Y(\reg_file_next[20][20] )
         );
  MXI2XL U954 ( .A(n1606), .B(n2180), .S0(n2983), .Y(\reg_file_next[16][20] )
         );
  MXI2XL U955 ( .A(n166), .B(n2180), .S0(n2970), .Y(\reg_file_next[28][20] )
         );
  MXI2XL U956 ( .A(n1991), .B(n2178), .S0(n2964), .Y(\reg_file_next[4][21] )
         );
  MXI2XL U957 ( .A(n2119), .B(n2178), .S0(n2990), .Y(\reg_file_next[0][21] )
         );
  MXI2XL U958 ( .A(n1735), .B(n2178), .S0(n2987), .Y(\reg_file_next[12][21] )
         );
  MXI2XL U959 ( .A(n1863), .B(n2178), .S0(n2960), .Y(\reg_file_next[8][21] )
         );
  MXI2XL U960 ( .A(n1479), .B(n2178), .S0(n2978), .Y(\reg_file_next[20][21] )
         );
  MXI2XL U961 ( .A(n1607), .B(n2178), .S0(n2983), .Y(\reg_file_next[16][21] )
         );
  MXI2XL U962 ( .A(n167), .B(n2178), .S0(n2970), .Y(\reg_file_next[28][21] )
         );
  MXI2XL U963 ( .A(n1992), .B(n2176), .S0(n2964), .Y(\reg_file_next[4][22] )
         );
  MXI2XL U964 ( .A(n2120), .B(n2176), .S0(n2990), .Y(\reg_file_next[0][22] )
         );
  MXI2XL U965 ( .A(n1736), .B(n2176), .S0(n2987), .Y(\reg_file_next[12][22] )
         );
  MXI2XL U966 ( .A(n1864), .B(n2176), .S0(n2960), .Y(\reg_file_next[8][22] )
         );
  MXI2XL U967 ( .A(n1480), .B(n2176), .S0(n2978), .Y(\reg_file_next[20][22] )
         );
  MXI2XL U968 ( .A(n1608), .B(n2176), .S0(n2983), .Y(\reg_file_next[16][22] )
         );
  MXI2XL U969 ( .A(n168), .B(n2176), .S0(n2970), .Y(\reg_file_next[28][22] )
         );
  MXI2XL U970 ( .A(n1993), .B(n2174), .S0(n2964), .Y(\reg_file_next[4][23] )
         );
  MXI2XL U971 ( .A(n2121), .B(n2174), .S0(n2990), .Y(\reg_file_next[0][23] )
         );
  MXI2XL U972 ( .A(n1737), .B(n2174), .S0(n2987), .Y(\reg_file_next[12][23] )
         );
  MXI2XL U973 ( .A(n1865), .B(n2174), .S0(n2960), .Y(\reg_file_next[8][23] )
         );
  MXI2XL U974 ( .A(n1481), .B(n2174), .S0(n2978), .Y(\reg_file_next[20][23] )
         );
  MXI2XL U975 ( .A(n1609), .B(n2174), .S0(n2983), .Y(\reg_file_next[16][23] )
         );
  MXI2XL U976 ( .A(n169), .B(n2174), .S0(n2970), .Y(\reg_file_next[28][23] )
         );
  MXI2XL U977 ( .A(n1994), .B(n2172), .S0(n2964), .Y(\reg_file_next[4][24] )
         );
  MXI2XL U978 ( .A(n2122), .B(n2172), .S0(n2990), .Y(\reg_file_next[0][24] )
         );
  MXI2XL U979 ( .A(n1738), .B(n2172), .S0(n2987), .Y(\reg_file_next[12][24] )
         );
  MXI2XL U980 ( .A(n1866), .B(n2172), .S0(n2960), .Y(\reg_file_next[8][24] )
         );
  MXI2XL U981 ( .A(n1482), .B(n2172), .S0(n2978), .Y(\reg_file_next[20][24] )
         );
  MXI2XL U982 ( .A(n1610), .B(n2172), .S0(n2983), .Y(\reg_file_next[16][24] )
         );
  MXI2XL U983 ( .A(n170), .B(n2172), .S0(n2970), .Y(\reg_file_next[28][24] )
         );
  MXI2XL U984 ( .A(n1995), .B(n2170), .S0(n2964), .Y(\reg_file_next[4][25] )
         );
  MXI2XL U985 ( .A(n2123), .B(n2170), .S0(n2990), .Y(\reg_file_next[0][25] )
         );
  MXI2XL U986 ( .A(n1739), .B(n2170), .S0(n2987), .Y(\reg_file_next[12][25] )
         );
  MXI2XL U987 ( .A(n1867), .B(n2170), .S0(n2960), .Y(\reg_file_next[8][25] )
         );
  MXI2XL U988 ( .A(n1483), .B(n2170), .S0(n2978), .Y(\reg_file_next[20][25] )
         );
  MXI2XL U989 ( .A(n1611), .B(n2170), .S0(n2983), .Y(\reg_file_next[16][25] )
         );
  MXI2XL U990 ( .A(n171), .B(n2170), .S0(n2970), .Y(\reg_file_next[28][25] )
         );
  MXI2XL U991 ( .A(n1996), .B(n2168), .S0(n2964), .Y(\reg_file_next[4][26] )
         );
  MXI2XL U992 ( .A(n2124), .B(n2168), .S0(n2990), .Y(\reg_file_next[0][26] )
         );
  MXI2XL U993 ( .A(n1740), .B(n2168), .S0(n2987), .Y(\reg_file_next[12][26] )
         );
  MXI2XL U994 ( .A(n1868), .B(n2168), .S0(n2960), .Y(\reg_file_next[8][26] )
         );
  MXI2XL U995 ( .A(n1484), .B(n2168), .S0(n2978), .Y(\reg_file_next[20][26] )
         );
  MXI2XL U996 ( .A(n1612), .B(n2168), .S0(n2983), .Y(\reg_file_next[16][26] )
         );
  MXI2XL U997 ( .A(n172), .B(n2168), .S0(n2970), .Y(\reg_file_next[28][26] )
         );
  MXI2XL U998 ( .A(n1997), .B(n2166), .S0(n2964), .Y(\reg_file_next[4][27] )
         );
  MXI2XL U999 ( .A(n2125), .B(n2166), .S0(n2990), .Y(\reg_file_next[0][27] )
         );
  MXI2XL U1000 ( .A(n1741), .B(n2166), .S0(n2987), .Y(\reg_file_next[12][27] )
         );
  MXI2XL U1001 ( .A(n1869), .B(n2166), .S0(n2960), .Y(\reg_file_next[8][27] )
         );
  MXI2XL U1002 ( .A(n1485), .B(n2166), .S0(n2978), .Y(\reg_file_next[20][27] )
         );
  MXI2XL U1003 ( .A(n1613), .B(n2166), .S0(n2983), .Y(\reg_file_next[16][27] )
         );
  MXI2XL U1004 ( .A(n173), .B(n2166), .S0(n2970), .Y(\reg_file_next[28][27] )
         );
  MXI2XL U1005 ( .A(n1998), .B(n2164), .S0(n2964), .Y(\reg_file_next[4][28] )
         );
  MXI2XL U1006 ( .A(n2126), .B(n2164), .S0(n2990), .Y(\reg_file_next[0][28] )
         );
  MXI2XL U1007 ( .A(n1742), .B(n2164), .S0(n2987), .Y(\reg_file_next[12][28] )
         );
  MXI2XL U1008 ( .A(n1870), .B(n2164), .S0(n2960), .Y(\reg_file_next[8][28] )
         );
  MXI2XL U1009 ( .A(n1486), .B(n2164), .S0(n2978), .Y(\reg_file_next[20][28] )
         );
  MXI2XL U1010 ( .A(n1614), .B(n2164), .S0(n2983), .Y(\reg_file_next[16][28] )
         );
  MXI2XL U1011 ( .A(n174), .B(n2164), .S0(n2970), .Y(\reg_file_next[28][28] )
         );
  MXI2XL U1012 ( .A(n1999), .B(n2162), .S0(n2964), .Y(\reg_file_next[4][29] )
         );
  MXI2XL U1013 ( .A(n2127), .B(n2162), .S0(n2990), .Y(\reg_file_next[0][29] )
         );
  MXI2XL U1014 ( .A(n1743), .B(n2162), .S0(n2987), .Y(\reg_file_next[12][29] )
         );
  MXI2XL U1015 ( .A(n1871), .B(n2162), .S0(n2960), .Y(\reg_file_next[8][29] )
         );
  MXI2XL U1016 ( .A(n1487), .B(n2162), .S0(n2978), .Y(\reg_file_next[20][29] )
         );
  MXI2XL U1017 ( .A(n1615), .B(n2162), .S0(n2983), .Y(\reg_file_next[16][29] )
         );
  MXI2XL U1018 ( .A(n175), .B(n2162), .S0(n2970), .Y(\reg_file_next[28][29] )
         );
  MXI2XL U1019 ( .A(n2000), .B(n2158), .S0(n2964), .Y(\reg_file_next[4][30] )
         );
  MXI2XL U1020 ( .A(n2128), .B(n2158), .S0(n2990), .Y(\reg_file_next[0][30] )
         );
  MXI2XL U1021 ( .A(n1744), .B(n2158), .S0(n2987), .Y(\reg_file_next[12][30] )
         );
  MXI2XL U1022 ( .A(n1872), .B(n2158), .S0(n2960), .Y(\reg_file_next[8][30] )
         );
  MXI2XL U1023 ( .A(n1488), .B(n2158), .S0(n2978), .Y(\reg_file_next[20][30] )
         );
  MXI2XL U1024 ( .A(n1616), .B(n2158), .S0(n2983), .Y(\reg_file_next[16][30] )
         );
  MXI2XL U1025 ( .A(n176), .B(n2158), .S0(n2970), .Y(\reg_file_next[28][30] )
         );
  MXI2XL U1026 ( .A(n2001), .B(n2156), .S0(n2964), .Y(\reg_file_next[4][31] )
         );
  MXI2XL U1027 ( .A(n2129), .B(n2156), .S0(n2990), .Y(\reg_file_next[0][31] )
         );
  MXI2XL U1028 ( .A(n1745), .B(n2156), .S0(n2987), .Y(\reg_file_next[12][31] )
         );
  MXI2XL U1029 ( .A(n1873), .B(n2156), .S0(n2960), .Y(\reg_file_next[8][31] )
         );
  MXI2XL U1030 ( .A(n1489), .B(n2156), .S0(n2978), .Y(\reg_file_next[20][31] )
         );
  MXI2XL U1031 ( .A(n1617), .B(n2156), .S0(n2983), .Y(\reg_file_next[16][31] )
         );
  MXI2XL U1032 ( .A(n177), .B(n2156), .S0(n2970), .Y(\reg_file_next[28][31] )
         );
  MXI2XL U1033 ( .A(n274), .B(n2204), .S0(n2974), .Y(\reg_file_next[24][0] )
         );
  MXI2XL U1034 ( .A(n275), .B(n2182), .S0(n2974), .Y(\reg_file_next[24][1] )
         );
  MXI2XL U1035 ( .A(n276), .B(n2160), .S0(n2974), .Y(\reg_file_next[24][2] )
         );
  MXI2XL U1036 ( .A(n277), .B(n2154), .S0(n2974), .Y(\reg_file_next[24][3] )
         );
  MXI2XL U1037 ( .A(n278), .B(n2152), .S0(n2974), .Y(\reg_file_next[24][4] )
         );
  MXI2XL U1038 ( .A(n279), .B(n2150), .S0(n2974), .Y(\reg_file_next[24][5] )
         );
  MXI2XL U1039 ( .A(n280), .B(n2148), .S0(n2974), .Y(\reg_file_next[24][6] )
         );
  MXI2XL U1040 ( .A(n281), .B(n2146), .S0(n2974), .Y(\reg_file_next[24][7] )
         );
  MXI2XL U1041 ( .A(n282), .B(n2144), .S0(n2974), .Y(\reg_file_next[24][8] )
         );
  MXI2XL U1042 ( .A(n283), .B(n2142), .S0(n2974), .Y(\reg_file_next[24][9] )
         );
  MXI2XL U1043 ( .A(n284), .B(n2202), .S0(n2974), .Y(\reg_file_next[24][10] )
         );
  MXI2XL U1044 ( .A(n285), .B(n2200), .S0(n2974), .Y(\reg_file_next[24][11] )
         );
  MXI2XL U1045 ( .A(n286), .B(n2198), .S0(n2974), .Y(\reg_file_next[24][12] )
         );
  MXI2XL U1046 ( .A(n287), .B(n2196), .S0(n2974), .Y(\reg_file_next[24][13] )
         );
  MXI2XL U1047 ( .A(n288), .B(n2194), .S0(n2974), .Y(\reg_file_next[24][14] )
         );
  MXI2XL U1048 ( .A(n289), .B(n2192), .S0(n2974), .Y(\reg_file_next[24][15] )
         );
  MXI2XL U1049 ( .A(n290), .B(n2190), .S0(n2974), .Y(\reg_file_next[24][16] )
         );
  MXI2XL U1050 ( .A(n291), .B(n2188), .S0(n2974), .Y(\reg_file_next[24][17] )
         );
  MXI2XL U1051 ( .A(n292), .B(n2186), .S0(n2974), .Y(\reg_file_next[24][18] )
         );
  MXI2XL U1052 ( .A(n293), .B(n2184), .S0(n2974), .Y(\reg_file_next[24][19] )
         );
  MXI2XL U1053 ( .A(n294), .B(n2180), .S0(n2974), .Y(\reg_file_next[24][20] )
         );
  MXI2XL U1054 ( .A(n295), .B(n2178), .S0(n2974), .Y(\reg_file_next[24][21] )
         );
  MXI2XL U1055 ( .A(n296), .B(n2176), .S0(n2974), .Y(\reg_file_next[24][22] )
         );
  MXI2XL U1056 ( .A(n297), .B(n2174), .S0(n2974), .Y(\reg_file_next[24][23] )
         );
  MXI2XL U1057 ( .A(n298), .B(n2172), .S0(n2974), .Y(\reg_file_next[24][24] )
         );
  MXI2XL U1058 ( .A(n1355), .B(n2170), .S0(n2974), .Y(\reg_file_next[24][25] )
         );
  MXI2XL U1059 ( .A(n1356), .B(n2168), .S0(n2974), .Y(\reg_file_next[24][26] )
         );
  MXI2XL U1060 ( .A(n1357), .B(n2166), .S0(n2974), .Y(\reg_file_next[24][27] )
         );
  MXI2XL U1061 ( .A(n1358), .B(n2164), .S0(n2974), .Y(\reg_file_next[24][28] )
         );
  MXI2XL U1062 ( .A(n1359), .B(n2162), .S0(n2974), .Y(\reg_file_next[24][29] )
         );
  MXI2XL U1063 ( .A(n1360), .B(n2158), .S0(n2974), .Y(\reg_file_next[24][30] )
         );
  MXI2XL U1064 ( .A(n1361), .B(n2156), .S0(n2974), .Y(\reg_file_next[24][31] )
         );
  MXI2XL U1065 ( .A(n1938), .B(n2204), .S0(n2963), .Y(\reg_file_next[5][0] )
         );
  MXI2XL U1066 ( .A(n2066), .B(n2204), .S0(n2979), .Y(\reg_file_next[1][0] )
         );
  MXI2XL U1067 ( .A(n1682), .B(n2204), .S0(n2986), .Y(\reg_file_next[13][0] )
         );
  MXI2XL U1068 ( .A(n1810), .B(n2204), .S0(n2928), .Y(\reg_file_next[9][0] )
         );
  MXI2XL U1069 ( .A(n1426), .B(n2204), .S0(n2977), .Y(\reg_file_next[21][0] )
         );
  MXI2XL U1070 ( .A(n1554), .B(n2204), .S0(n2982), .Y(\reg_file_next[17][0] )
         );
  MXI2XL U1071 ( .A(n114), .B(n2204), .S0(n2969), .Y(\reg_file_next[29][0] )
         );
  MXI2XL U1072 ( .A(n1939), .B(n2182), .S0(n2963), .Y(\reg_file_next[5][1] )
         );
  MXI2XL U1073 ( .A(n2067), .B(n2182), .S0(n2979), .Y(\reg_file_next[1][1] )
         );
  MXI2XL U1074 ( .A(n1683), .B(n2182), .S0(n2986), .Y(\reg_file_next[13][1] )
         );
  MXI2XL U1075 ( .A(n1811), .B(n2182), .S0(n2928), .Y(\reg_file_next[9][1] )
         );
  MXI2XL U1076 ( .A(n1427), .B(n2182), .S0(n2977), .Y(\reg_file_next[21][1] )
         );
  MXI2XL U1077 ( .A(n1555), .B(n2182), .S0(n2982), .Y(\reg_file_next[17][1] )
         );
  MXI2XL U1078 ( .A(n115), .B(n2182), .S0(n2969), .Y(\reg_file_next[29][1] )
         );
  MXI2XL U1079 ( .A(n1940), .B(n2160), .S0(n2963), .Y(\reg_file_next[5][2] )
         );
  MXI2XL U1080 ( .A(n2068), .B(n2160), .S0(n2979), .Y(\reg_file_next[1][2] )
         );
  MXI2XL U1081 ( .A(n1684), .B(n2160), .S0(n2986), .Y(\reg_file_next[13][2] )
         );
  MXI2XL U1082 ( .A(n1812), .B(n2160), .S0(n2928), .Y(\reg_file_next[9][2] )
         );
  MXI2XL U1083 ( .A(n1428), .B(n2160), .S0(n2977), .Y(\reg_file_next[21][2] )
         );
  MXI2XL U1084 ( .A(n1556), .B(n2160), .S0(n2982), .Y(\reg_file_next[17][2] )
         );
  MXI2XL U1085 ( .A(n116), .B(n2160), .S0(n2969), .Y(\reg_file_next[29][2] )
         );
  MXI2XL U1086 ( .A(n1941), .B(n2154), .S0(n2963), .Y(\reg_file_next[5][3] )
         );
  MXI2XL U1087 ( .A(n2069), .B(n2154), .S0(n2979), .Y(\reg_file_next[1][3] )
         );
  MXI2XL U1088 ( .A(n1685), .B(n2154), .S0(n2986), .Y(\reg_file_next[13][3] )
         );
  MXI2XL U1089 ( .A(n1813), .B(n2154), .S0(n2928), .Y(\reg_file_next[9][3] )
         );
  MXI2XL U1090 ( .A(n1429), .B(n2154), .S0(n2977), .Y(\reg_file_next[21][3] )
         );
  MXI2XL U1091 ( .A(n1557), .B(n2154), .S0(n2982), .Y(\reg_file_next[17][3] )
         );
  MXI2XL U1092 ( .A(n117), .B(n2154), .S0(n2969), .Y(\reg_file_next[29][3] )
         );
  MXI2XL U1093 ( .A(n1942), .B(n2152), .S0(n2963), .Y(\reg_file_next[5][4] )
         );
  MXI2XL U1094 ( .A(n2070), .B(n2152), .S0(n2979), .Y(\reg_file_next[1][4] )
         );
  MXI2XL U1095 ( .A(n1686), .B(n2152), .S0(n2986), .Y(\reg_file_next[13][4] )
         );
  MXI2XL U1096 ( .A(n1814), .B(n2152), .S0(n2928), .Y(\reg_file_next[9][4] )
         );
  MXI2XL U1097 ( .A(n1430), .B(n2152), .S0(n2977), .Y(\reg_file_next[21][4] )
         );
  MXI2XL U1098 ( .A(n1558), .B(n2152), .S0(n2982), .Y(\reg_file_next[17][4] )
         );
  MXI2XL U1099 ( .A(n118), .B(n2152), .S0(n2969), .Y(\reg_file_next[29][4] )
         );
  MXI2XL U1100 ( .A(n1943), .B(n2150), .S0(n2963), .Y(\reg_file_next[5][5] )
         );
  MXI2XL U1101 ( .A(n2071), .B(n2150), .S0(n2979), .Y(\reg_file_next[1][5] )
         );
  MXI2XL U1102 ( .A(n1687), .B(n2150), .S0(n2986), .Y(\reg_file_next[13][5] )
         );
  MXI2XL U1103 ( .A(n1815), .B(n2150), .S0(n2928), .Y(\reg_file_next[9][5] )
         );
  MXI2XL U1104 ( .A(n1431), .B(n2150), .S0(n2977), .Y(\reg_file_next[21][5] )
         );
  MXI2XL U1105 ( .A(n1559), .B(n2150), .S0(n2982), .Y(\reg_file_next[17][5] )
         );
  MXI2XL U1106 ( .A(n119), .B(n2150), .S0(n2969), .Y(\reg_file_next[29][5] )
         );
  MXI2XL U1107 ( .A(n1944), .B(n2148), .S0(n2963), .Y(\reg_file_next[5][6] )
         );
  MXI2XL U1108 ( .A(n2072), .B(n2148), .S0(n2979), .Y(\reg_file_next[1][6] )
         );
  MXI2XL U1109 ( .A(n1688), .B(n2148), .S0(n2986), .Y(\reg_file_next[13][6] )
         );
  MXI2XL U1110 ( .A(n1816), .B(n2148), .S0(n2928), .Y(\reg_file_next[9][6] )
         );
  MXI2XL U1111 ( .A(n1432), .B(n2148), .S0(n2977), .Y(\reg_file_next[21][6] )
         );
  MXI2XL U1112 ( .A(n1560), .B(n2148), .S0(n2982), .Y(\reg_file_next[17][6] )
         );
  MXI2XL U1113 ( .A(n120), .B(n2148), .S0(n2969), .Y(\reg_file_next[29][6] )
         );
  MXI2XL U1114 ( .A(n1945), .B(n2146), .S0(n2963), .Y(\reg_file_next[5][7] )
         );
  MXI2XL U1115 ( .A(n2073), .B(n2146), .S0(n2979), .Y(\reg_file_next[1][7] )
         );
  MXI2XL U1116 ( .A(n1689), .B(n2146), .S0(n2986), .Y(\reg_file_next[13][7] )
         );
  MXI2XL U1117 ( .A(n1817), .B(n2146), .S0(n2928), .Y(\reg_file_next[9][7] )
         );
  MXI2XL U1118 ( .A(n1433), .B(n2146), .S0(n2977), .Y(\reg_file_next[21][7] )
         );
  MXI2XL U1119 ( .A(n1561), .B(n2146), .S0(n2982), .Y(\reg_file_next[17][7] )
         );
  MXI2XL U1120 ( .A(n121), .B(n2146), .S0(n2969), .Y(\reg_file_next[29][7] )
         );
  MXI2XL U1121 ( .A(n1946), .B(n2144), .S0(n2963), .Y(\reg_file_next[5][8] )
         );
  MXI2XL U1122 ( .A(n2074), .B(n2144), .S0(n2979), .Y(\reg_file_next[1][8] )
         );
  MXI2XL U1123 ( .A(n1690), .B(n2144), .S0(n2986), .Y(\reg_file_next[13][8] )
         );
  MXI2XL U1124 ( .A(n1818), .B(n2144), .S0(n2928), .Y(\reg_file_next[9][8] )
         );
  MXI2XL U1125 ( .A(n1434), .B(n2144), .S0(n2977), .Y(\reg_file_next[21][8] )
         );
  MXI2XL U1126 ( .A(n1562), .B(n2144), .S0(n2982), .Y(\reg_file_next[17][8] )
         );
  MXI2XL U1127 ( .A(n122), .B(n2144), .S0(n2969), .Y(\reg_file_next[29][8] )
         );
  MXI2XL U1128 ( .A(n1947), .B(n2142), .S0(n2963), .Y(\reg_file_next[5][9] )
         );
  MXI2XL U1129 ( .A(n2075), .B(n2142), .S0(n2979), .Y(\reg_file_next[1][9] )
         );
  MXI2XL U1130 ( .A(n1691), .B(n2142), .S0(n2986), .Y(\reg_file_next[13][9] )
         );
  MXI2XL U1131 ( .A(n1819), .B(n2142), .S0(n2928), .Y(\reg_file_next[9][9] )
         );
  MXI2XL U1132 ( .A(n1435), .B(n2142), .S0(n2977), .Y(\reg_file_next[21][9] )
         );
  MXI2XL U1133 ( .A(n1563), .B(n2142), .S0(n2982), .Y(\reg_file_next[17][9] )
         );
  MXI2XL U1134 ( .A(n123), .B(n2142), .S0(n2969), .Y(\reg_file_next[29][9] )
         );
  MXI2XL U1135 ( .A(n1948), .B(n2202), .S0(n2963), .Y(\reg_file_next[5][10] )
         );
  MXI2XL U1136 ( .A(n2076), .B(n2202), .S0(n2979), .Y(\reg_file_next[1][10] )
         );
  MXI2XL U1137 ( .A(n1692), .B(n2202), .S0(n2986), .Y(\reg_file_next[13][10] )
         );
  MXI2XL U1138 ( .A(n1820), .B(n2202), .S0(n2928), .Y(\reg_file_next[9][10] )
         );
  MXI2XL U1139 ( .A(n1436), .B(n2202), .S0(n2977), .Y(\reg_file_next[21][10] )
         );
  MXI2XL U1140 ( .A(n1564), .B(n2202), .S0(n2982), .Y(\reg_file_next[17][10] )
         );
  MXI2XL U1141 ( .A(n124), .B(n2202), .S0(n2969), .Y(\reg_file_next[29][10] )
         );
  MXI2XL U1142 ( .A(n1949), .B(n2200), .S0(n2963), .Y(\reg_file_next[5][11] )
         );
  MXI2XL U1143 ( .A(n2077), .B(n2200), .S0(n2979), .Y(\reg_file_next[1][11] )
         );
  MXI2XL U1144 ( .A(n1693), .B(n2200), .S0(n2986), .Y(\reg_file_next[13][11] )
         );
  MXI2XL U1145 ( .A(n1821), .B(n2200), .S0(n2928), .Y(\reg_file_next[9][11] )
         );
  MXI2XL U1146 ( .A(n1437), .B(n2200), .S0(n2977), .Y(\reg_file_next[21][11] )
         );
  MXI2XL U1147 ( .A(n1565), .B(n2200), .S0(n2982), .Y(\reg_file_next[17][11] )
         );
  MXI2XL U1148 ( .A(n125), .B(n2200), .S0(n2969), .Y(\reg_file_next[29][11] )
         );
  MXI2XL U1149 ( .A(n1950), .B(n2198), .S0(n2963), .Y(\reg_file_next[5][12] )
         );
  MXI2XL U1150 ( .A(n2078), .B(n2198), .S0(n2979), .Y(\reg_file_next[1][12] )
         );
  MXI2XL U1151 ( .A(n1694), .B(n2198), .S0(n2986), .Y(\reg_file_next[13][12] )
         );
  MXI2XL U1152 ( .A(n1822), .B(n2198), .S0(n2928), .Y(\reg_file_next[9][12] )
         );
  MXI2XL U1153 ( .A(n1438), .B(n2198), .S0(n2977), .Y(\reg_file_next[21][12] )
         );
  MXI2XL U1154 ( .A(n1566), .B(n2198), .S0(n2982), .Y(\reg_file_next[17][12] )
         );
  MXI2XL U1155 ( .A(n126), .B(n2198), .S0(n2969), .Y(\reg_file_next[29][12] )
         );
  MXI2XL U1156 ( .A(n1951), .B(n2196), .S0(n2963), .Y(\reg_file_next[5][13] )
         );
  MXI2XL U1157 ( .A(n2079), .B(n2196), .S0(n2979), .Y(\reg_file_next[1][13] )
         );
  MXI2XL U1158 ( .A(n1695), .B(n2196), .S0(n2986), .Y(\reg_file_next[13][13] )
         );
  MXI2XL U1159 ( .A(n1823), .B(n2196), .S0(n2928), .Y(\reg_file_next[9][13] )
         );
  MXI2XL U1160 ( .A(n1439), .B(n2196), .S0(n2977), .Y(\reg_file_next[21][13] )
         );
  MXI2XL U1161 ( .A(n1567), .B(n2196), .S0(n2982), .Y(\reg_file_next[17][13] )
         );
  MXI2XL U1162 ( .A(n127), .B(n2196), .S0(n2969), .Y(\reg_file_next[29][13] )
         );
  MXI2XL U1163 ( .A(n1952), .B(n2194), .S0(n2963), .Y(\reg_file_next[5][14] )
         );
  MXI2XL U1164 ( .A(n2080), .B(n2194), .S0(n2979), .Y(\reg_file_next[1][14] )
         );
  MXI2XL U1165 ( .A(n1696), .B(n2194), .S0(n2986), .Y(\reg_file_next[13][14] )
         );
  MXI2XL U1166 ( .A(n1824), .B(n2194), .S0(n2928), .Y(\reg_file_next[9][14] )
         );
  MXI2XL U1167 ( .A(n1440), .B(n2194), .S0(n2977), .Y(\reg_file_next[21][14] )
         );
  MXI2XL U1168 ( .A(n1568), .B(n2194), .S0(n2982), .Y(\reg_file_next[17][14] )
         );
  MXI2XL U1169 ( .A(n128), .B(n2194), .S0(n2969), .Y(\reg_file_next[29][14] )
         );
  MXI2XL U1170 ( .A(n1953), .B(n2192), .S0(n2963), .Y(\reg_file_next[5][15] )
         );
  MXI2XL U1171 ( .A(n2081), .B(n2192), .S0(n2979), .Y(\reg_file_next[1][15] )
         );
  MXI2XL U1172 ( .A(n1697), .B(n2192), .S0(n2986), .Y(\reg_file_next[13][15] )
         );
  MXI2XL U1173 ( .A(n1825), .B(n2192), .S0(n2928), .Y(\reg_file_next[9][15] )
         );
  MXI2XL U1174 ( .A(n1441), .B(n2192), .S0(n2977), .Y(\reg_file_next[21][15] )
         );
  MXI2XL U1175 ( .A(n1569), .B(n2192), .S0(n2982), .Y(\reg_file_next[17][15] )
         );
  MXI2XL U1176 ( .A(n129), .B(n2192), .S0(n2969), .Y(\reg_file_next[29][15] )
         );
  MXI2XL U1177 ( .A(n1954), .B(n2190), .S0(n2963), .Y(\reg_file_next[5][16] )
         );
  MXI2XL U1178 ( .A(n2082), .B(n2190), .S0(n2979), .Y(\reg_file_next[1][16] )
         );
  MXI2XL U1179 ( .A(n1698), .B(n2190), .S0(n2986), .Y(\reg_file_next[13][16] )
         );
  MXI2XL U1180 ( .A(n1826), .B(n2190), .S0(n2928), .Y(\reg_file_next[9][16] )
         );
  MXI2XL U1181 ( .A(n1442), .B(n2190), .S0(n2977), .Y(\reg_file_next[21][16] )
         );
  MXI2XL U1182 ( .A(n1570), .B(n2190), .S0(n2982), .Y(\reg_file_next[17][16] )
         );
  MXI2XL U1183 ( .A(n130), .B(n2190), .S0(n2969), .Y(\reg_file_next[29][16] )
         );
  MXI2XL U1184 ( .A(n1955), .B(n2188), .S0(n2963), .Y(\reg_file_next[5][17] )
         );
  MXI2XL U1185 ( .A(n2083), .B(n2188), .S0(n2979), .Y(\reg_file_next[1][17] )
         );
  MXI2XL U1186 ( .A(n1699), .B(n2188), .S0(n2986), .Y(\reg_file_next[13][17] )
         );
  MXI2XL U1187 ( .A(n1827), .B(n2188), .S0(n2928), .Y(\reg_file_next[9][17] )
         );
  MXI2XL U1188 ( .A(n1443), .B(n2188), .S0(n2977), .Y(\reg_file_next[21][17] )
         );
  MXI2XL U1189 ( .A(n1571), .B(n2188), .S0(n2982), .Y(\reg_file_next[17][17] )
         );
  MXI2XL U1190 ( .A(n131), .B(n2188), .S0(n2969), .Y(\reg_file_next[29][17] )
         );
  MXI2XL U1191 ( .A(n1956), .B(n2186), .S0(n2963), .Y(\reg_file_next[5][18] )
         );
  MXI2XL U1192 ( .A(n2084), .B(n2186), .S0(n2979), .Y(\reg_file_next[1][18] )
         );
  MXI2XL U1193 ( .A(n1700), .B(n2186), .S0(n2986), .Y(\reg_file_next[13][18] )
         );
  MXI2XL U1194 ( .A(n1828), .B(n2186), .S0(n2928), .Y(\reg_file_next[9][18] )
         );
  MXI2XL U1195 ( .A(n1444), .B(n2186), .S0(n2977), .Y(\reg_file_next[21][18] )
         );
  MXI2XL U1196 ( .A(n1572), .B(n2186), .S0(n2982), .Y(\reg_file_next[17][18] )
         );
  MXI2XL U1197 ( .A(n132), .B(n2186), .S0(n2969), .Y(\reg_file_next[29][18] )
         );
  MXI2XL U1198 ( .A(n1957), .B(n2184), .S0(n2963), .Y(\reg_file_next[5][19] )
         );
  MXI2XL U1199 ( .A(n2085), .B(n2184), .S0(n2979), .Y(\reg_file_next[1][19] )
         );
  MXI2XL U1200 ( .A(n1701), .B(n2184), .S0(n2986), .Y(\reg_file_next[13][19] )
         );
  MXI2XL U1201 ( .A(n1829), .B(n2184), .S0(n2928), .Y(\reg_file_next[9][19] )
         );
  MXI2XL U1202 ( .A(n1445), .B(n2184), .S0(n2977), .Y(\reg_file_next[21][19] )
         );
  MXI2XL U1203 ( .A(n1573), .B(n2184), .S0(n2982), .Y(\reg_file_next[17][19] )
         );
  MXI2XL U1204 ( .A(n133), .B(n2184), .S0(n2969), .Y(\reg_file_next[29][19] )
         );
  MXI2XL U1205 ( .A(n1958), .B(n2180), .S0(n2963), .Y(\reg_file_next[5][20] )
         );
  MXI2XL U1206 ( .A(n2086), .B(n2180), .S0(n2979), .Y(\reg_file_next[1][20] )
         );
  MXI2XL U1207 ( .A(n1702), .B(n2180), .S0(n2986), .Y(\reg_file_next[13][20] )
         );
  MXI2XL U1208 ( .A(n1830), .B(n2180), .S0(n2928), .Y(\reg_file_next[9][20] )
         );
  MXI2XL U1209 ( .A(n1446), .B(n2180), .S0(n2977), .Y(\reg_file_next[21][20] )
         );
  MXI2XL U1210 ( .A(n1574), .B(n2180), .S0(n2982), .Y(\reg_file_next[17][20] )
         );
  MXI2XL U1211 ( .A(n134), .B(n2180), .S0(n2969), .Y(\reg_file_next[29][20] )
         );
  MXI2XL U1212 ( .A(n1959), .B(n2178), .S0(n2963), .Y(\reg_file_next[5][21] )
         );
  MXI2XL U1213 ( .A(n2087), .B(n2178), .S0(n2979), .Y(\reg_file_next[1][21] )
         );
  MXI2XL U1214 ( .A(n1703), .B(n2178), .S0(n2986), .Y(\reg_file_next[13][21] )
         );
  MXI2XL U1215 ( .A(n1831), .B(n2178), .S0(n2928), .Y(\reg_file_next[9][21] )
         );
  MXI2XL U1216 ( .A(n1447), .B(n2178), .S0(n2977), .Y(\reg_file_next[21][21] )
         );
  MXI2XL U1217 ( .A(n1575), .B(n2178), .S0(n2982), .Y(\reg_file_next[17][21] )
         );
  MXI2XL U1218 ( .A(n135), .B(n2178), .S0(n2969), .Y(\reg_file_next[29][21] )
         );
  MXI2XL U1219 ( .A(n1960), .B(n2176), .S0(n2963), .Y(\reg_file_next[5][22] )
         );
  MXI2XL U1220 ( .A(n2088), .B(n2176), .S0(n2979), .Y(\reg_file_next[1][22] )
         );
  MXI2XL U1221 ( .A(n1704), .B(n2176), .S0(n2986), .Y(\reg_file_next[13][22] )
         );
  MXI2XL U1222 ( .A(n1832), .B(n2176), .S0(n2928), .Y(\reg_file_next[9][22] )
         );
  MXI2XL U1223 ( .A(n1448), .B(n2176), .S0(n2977), .Y(\reg_file_next[21][22] )
         );
  MXI2XL U1224 ( .A(n1576), .B(n2176), .S0(n2982), .Y(\reg_file_next[17][22] )
         );
  MXI2XL U1225 ( .A(n136), .B(n2176), .S0(n2969), .Y(\reg_file_next[29][22] )
         );
  MXI2XL U1226 ( .A(n1961), .B(n2174), .S0(n2963), .Y(\reg_file_next[5][23] )
         );
  MXI2XL U1227 ( .A(n2089), .B(n2174), .S0(n2979), .Y(\reg_file_next[1][23] )
         );
  MXI2XL U1228 ( .A(n1705), .B(n2174), .S0(n2986), .Y(\reg_file_next[13][23] )
         );
  MXI2XL U1229 ( .A(n1833), .B(n2174), .S0(n2928), .Y(\reg_file_next[9][23] )
         );
  MXI2XL U1230 ( .A(n1449), .B(n2174), .S0(n2977), .Y(\reg_file_next[21][23] )
         );
  MXI2XL U1231 ( .A(n1577), .B(n2174), .S0(n2982), .Y(\reg_file_next[17][23] )
         );
  MXI2XL U1232 ( .A(n137), .B(n2174), .S0(n2969), .Y(\reg_file_next[29][23] )
         );
  MXI2XL U1233 ( .A(n1962), .B(n2172), .S0(n2963), .Y(\reg_file_next[5][24] )
         );
  MXI2XL U1234 ( .A(n2090), .B(n2172), .S0(n2979), .Y(\reg_file_next[1][24] )
         );
  MXI2XL U1235 ( .A(n1706), .B(n2172), .S0(n2986), .Y(\reg_file_next[13][24] )
         );
  MXI2XL U1236 ( .A(n1834), .B(n2172), .S0(n2928), .Y(\reg_file_next[9][24] )
         );
  MXI2XL U1237 ( .A(n1450), .B(n2172), .S0(n2977), .Y(\reg_file_next[21][24] )
         );
  MXI2XL U1238 ( .A(n1578), .B(n2172), .S0(n2982), .Y(\reg_file_next[17][24] )
         );
  MXI2XL U1239 ( .A(n138), .B(n2172), .S0(n2969), .Y(\reg_file_next[29][24] )
         );
  MXI2XL U1240 ( .A(n1963), .B(n2170), .S0(n2963), .Y(\reg_file_next[5][25] )
         );
  MXI2XL U1241 ( .A(n2091), .B(n2170), .S0(n2979), .Y(\reg_file_next[1][25] )
         );
  MXI2XL U1242 ( .A(n1707), .B(n2170), .S0(n2986), .Y(\reg_file_next[13][25] )
         );
  MXI2XL U1243 ( .A(n1835), .B(n2170), .S0(n2928), .Y(\reg_file_next[9][25] )
         );
  MXI2XL U1244 ( .A(n1451), .B(n2170), .S0(n2977), .Y(\reg_file_next[21][25] )
         );
  MXI2XL U1245 ( .A(n1579), .B(n2170), .S0(n2982), .Y(\reg_file_next[17][25] )
         );
  MXI2XL U1246 ( .A(n139), .B(n2170), .S0(n2969), .Y(\reg_file_next[29][25] )
         );
  MXI2XL U1247 ( .A(n1964), .B(n2168), .S0(n2963), .Y(\reg_file_next[5][26] )
         );
  MXI2XL U1248 ( .A(n2092), .B(n2168), .S0(n2979), .Y(\reg_file_next[1][26] )
         );
  MXI2XL U1249 ( .A(n1708), .B(n2168), .S0(n2986), .Y(\reg_file_next[13][26] )
         );
  MXI2XL U1250 ( .A(n1836), .B(n2168), .S0(n2928), .Y(\reg_file_next[9][26] )
         );
  MXI2XL U1251 ( .A(n1452), .B(n2168), .S0(n2977), .Y(\reg_file_next[21][26] )
         );
  MXI2XL U1252 ( .A(n1580), .B(n2168), .S0(n2982), .Y(\reg_file_next[17][26] )
         );
  MXI2XL U1253 ( .A(n140), .B(n2168), .S0(n2969), .Y(\reg_file_next[29][26] )
         );
  MXI2XL U1254 ( .A(n1965), .B(n2166), .S0(n2963), .Y(\reg_file_next[5][27] )
         );
  MXI2XL U1255 ( .A(n2093), .B(n2166), .S0(n2979), .Y(\reg_file_next[1][27] )
         );
  MXI2XL U1256 ( .A(n1709), .B(n2166), .S0(n2986), .Y(\reg_file_next[13][27] )
         );
  MXI2XL U1257 ( .A(n1837), .B(n2166), .S0(n2928), .Y(\reg_file_next[9][27] )
         );
  MXI2XL U1258 ( .A(n1453), .B(n2166), .S0(n2977), .Y(\reg_file_next[21][27] )
         );
  MXI2XL U1259 ( .A(n1581), .B(n2166), .S0(n2982), .Y(\reg_file_next[17][27] )
         );
  MXI2XL U1260 ( .A(n141), .B(n2166), .S0(n2969), .Y(\reg_file_next[29][27] )
         );
  MXI2XL U1261 ( .A(n1966), .B(n2164), .S0(n2963), .Y(\reg_file_next[5][28] )
         );
  MXI2XL U1262 ( .A(n2094), .B(n2164), .S0(n2979), .Y(\reg_file_next[1][28] )
         );
  MXI2XL U1263 ( .A(n1710), .B(n2164), .S0(n2986), .Y(\reg_file_next[13][28] )
         );
  MXI2XL U1264 ( .A(n1838), .B(n2164), .S0(n2928), .Y(\reg_file_next[9][28] )
         );
  MXI2XL U1265 ( .A(n1454), .B(n2164), .S0(n2977), .Y(\reg_file_next[21][28] )
         );
  MXI2XL U1266 ( .A(n1582), .B(n2164), .S0(n2982), .Y(\reg_file_next[17][28] )
         );
  MXI2XL U1267 ( .A(n142), .B(n2164), .S0(n2969), .Y(\reg_file_next[29][28] )
         );
  MXI2XL U1268 ( .A(n1967), .B(n2162), .S0(n2963), .Y(\reg_file_next[5][29] )
         );
  MXI2XL U1269 ( .A(n2095), .B(n2162), .S0(n2979), .Y(\reg_file_next[1][29] )
         );
  MXI2XL U1270 ( .A(n1711), .B(n2162), .S0(n2986), .Y(\reg_file_next[13][29] )
         );
  MXI2XL U1271 ( .A(n1839), .B(n2162), .S0(n2928), .Y(\reg_file_next[9][29] )
         );
  MXI2XL U1272 ( .A(n1455), .B(n2162), .S0(n2977), .Y(\reg_file_next[21][29] )
         );
  MXI2XL U1273 ( .A(n1583), .B(n2162), .S0(n2982), .Y(\reg_file_next[17][29] )
         );
  MXI2XL U1274 ( .A(n143), .B(n2162), .S0(n2969), .Y(\reg_file_next[29][29] )
         );
  MXI2XL U1275 ( .A(n1968), .B(n2158), .S0(n2963), .Y(\reg_file_next[5][30] )
         );
  MXI2XL U1276 ( .A(n2096), .B(n2158), .S0(n2979), .Y(\reg_file_next[1][30] )
         );
  MXI2XL U1277 ( .A(n1712), .B(n2158), .S0(n2986), .Y(\reg_file_next[13][30] )
         );
  MXI2XL U1278 ( .A(n1840), .B(n2158), .S0(n2928), .Y(\reg_file_next[9][30] )
         );
  MXI2XL U1279 ( .A(n1456), .B(n2158), .S0(n2977), .Y(\reg_file_next[21][30] )
         );
  MXI2XL U1280 ( .A(n1584), .B(n2158), .S0(n2982), .Y(\reg_file_next[17][30] )
         );
  MXI2XL U1281 ( .A(n144), .B(n2158), .S0(n2969), .Y(\reg_file_next[29][30] )
         );
  MXI2XL U1282 ( .A(n1969), .B(n2156), .S0(n2963), .Y(\reg_file_next[5][31] )
         );
  MXI2XL U1283 ( .A(n2097), .B(n2156), .S0(n2979), .Y(\reg_file_next[1][31] )
         );
  MXI2XL U1284 ( .A(n1713), .B(n2156), .S0(n2986), .Y(\reg_file_next[13][31] )
         );
  MXI2XL U1285 ( .A(n1841), .B(n2156), .S0(n2928), .Y(\reg_file_next[9][31] )
         );
  MXI2XL U1286 ( .A(n1457), .B(n2156), .S0(n2977), .Y(\reg_file_next[21][31] )
         );
  MXI2XL U1287 ( .A(n1585), .B(n2156), .S0(n2982), .Y(\reg_file_next[17][31] )
         );
  MXI2XL U1288 ( .A(n145), .B(n2156), .S0(n2969), .Y(\reg_file_next[29][31] )
         );
  MXI2XL U1289 ( .A(n242), .B(n2204), .S0(n2973), .Y(\reg_file_next[25][0] )
         );
  MXI2XL U1290 ( .A(n243), .B(n2182), .S0(n2973), .Y(\reg_file_next[25][1] )
         );
  MXI2XL U1291 ( .A(n244), .B(n2160), .S0(n2973), .Y(\reg_file_next[25][2] )
         );
  MXI2XL U1292 ( .A(n245), .B(n2154), .S0(n2973), .Y(\reg_file_next[25][3] )
         );
  MXI2XL U1293 ( .A(n246), .B(n2152), .S0(n2973), .Y(\reg_file_next[25][4] )
         );
  MXI2XL U1294 ( .A(n247), .B(n2150), .S0(n2973), .Y(\reg_file_next[25][5] )
         );
  MXI2XL U1295 ( .A(n248), .B(n2148), .S0(n2973), .Y(\reg_file_next[25][6] )
         );
  MXI2XL U1296 ( .A(n249), .B(n2146), .S0(n2973), .Y(\reg_file_next[25][7] )
         );
  MXI2XL U1297 ( .A(n250), .B(n2144), .S0(n2973), .Y(\reg_file_next[25][8] )
         );
  MXI2XL U1298 ( .A(n251), .B(n2142), .S0(n2973), .Y(\reg_file_next[25][9] )
         );
  MXI2XL U1299 ( .A(n252), .B(n2202), .S0(n2973), .Y(\reg_file_next[25][10] )
         );
  MXI2XL U1300 ( .A(n253), .B(n2200), .S0(n2973), .Y(\reg_file_next[25][11] )
         );
  MXI2XL U1301 ( .A(n254), .B(n2198), .S0(n2973), .Y(\reg_file_next[25][12] )
         );
  MXI2XL U1302 ( .A(n255), .B(n2196), .S0(n2973), .Y(\reg_file_next[25][13] )
         );
  MXI2XL U1303 ( .A(n256), .B(n2194), .S0(n2973), .Y(\reg_file_next[25][14] )
         );
  MXI2XL U1304 ( .A(n257), .B(n2192), .S0(n2973), .Y(\reg_file_next[25][15] )
         );
  MXI2XL U1305 ( .A(n258), .B(n2190), .S0(n2973), .Y(\reg_file_next[25][16] )
         );
  MXI2XL U1306 ( .A(n259), .B(n2188), .S0(n2973), .Y(\reg_file_next[25][17] )
         );
  MXI2XL U1307 ( .A(n260), .B(n2186), .S0(n2973), .Y(\reg_file_next[25][18] )
         );
  MXI2XL U1308 ( .A(n261), .B(n2184), .S0(n2973), .Y(\reg_file_next[25][19] )
         );
  MXI2XL U1309 ( .A(n262), .B(n2180), .S0(n2973), .Y(\reg_file_next[25][20] )
         );
  MXI2XL U1310 ( .A(n263), .B(n2178), .S0(n2973), .Y(\reg_file_next[25][21] )
         );
  MXI2XL U1311 ( .A(n264), .B(n2176), .S0(n2973), .Y(\reg_file_next[25][22] )
         );
  MXI2XL U1312 ( .A(n265), .B(n2174), .S0(n2973), .Y(\reg_file_next[25][23] )
         );
  MXI2XL U1313 ( .A(n266), .B(n2172), .S0(n2973), .Y(\reg_file_next[25][24] )
         );
  MXI2XL U1314 ( .A(n267), .B(n2170), .S0(n2973), .Y(\reg_file_next[25][25] )
         );
  MXI2XL U1315 ( .A(n268), .B(n2168), .S0(n2973), .Y(\reg_file_next[25][26] )
         );
  MXI2XL U1316 ( .A(n269), .B(n2166), .S0(n2973), .Y(\reg_file_next[25][27] )
         );
  MXI2XL U1317 ( .A(n270), .B(n2164), .S0(n2973), .Y(\reg_file_next[25][28] )
         );
  MXI2XL U1318 ( .A(n271), .B(n2162), .S0(n2973), .Y(\reg_file_next[25][29] )
         );
  MXI2XL U1319 ( .A(n272), .B(n2158), .S0(n2973), .Y(\reg_file_next[25][30] )
         );
  MXI2XL U1320 ( .A(n273), .B(n2156), .S0(n2973), .Y(\reg_file_next[25][31] )
         );
  NOR2BXL U1321 ( .AN(n2139), .B(Jump[1]), .Y(n3101) );
  MXI2XL U1322 ( .A(n49), .B(n2204), .S0(n3102), .Y(n1322) );
  MXI2XL U1323 ( .A(n50), .B(n2182), .S0(n3102), .Y(n1321) );
  MXI2XL U1324 ( .A(n51), .B(n2160), .S0(n3102), .Y(n1320) );
  MXI2XL U1325 ( .A(n52), .B(n2154), .S0(n3102), .Y(n1319) );
  MXI2XL U1326 ( .A(n53), .B(n2152), .S0(n3102), .Y(n1318) );
  MXI2XL U1327 ( .A(n54), .B(n2150), .S0(n3102), .Y(n1317) );
  MXI2XL U1328 ( .A(n55), .B(n2148), .S0(n3102), .Y(n1316) );
  MXI2XL U1329 ( .A(n56), .B(n2146), .S0(n3102), .Y(n1315) );
  MXI2XL U1330 ( .A(n57), .B(n2144), .S0(n3102), .Y(n1314) );
  MXI2XL U1331 ( .A(n58), .B(n2142), .S0(n3102), .Y(n1313) );
  MXI2XL U1332 ( .A(n59), .B(n2202), .S0(n3102), .Y(n1312) );
  MXI2XL U1333 ( .A(n60), .B(n2200), .S0(n3102), .Y(n1311) );
  MXI2XL U1334 ( .A(n61), .B(n2198), .S0(n3102), .Y(n1310) );
  MXI2XL U1335 ( .A(n62), .B(n2196), .S0(n3102), .Y(n1309) );
  MXI2XL U1336 ( .A(n63), .B(n2194), .S0(n3102), .Y(n1308) );
  MXI2XL U1337 ( .A(n64), .B(n2192), .S0(n3102), .Y(n1307) );
  MXI2XL U1338 ( .A(n65), .B(n2190), .S0(n3102), .Y(n1306) );
  MXI2XL U1339 ( .A(n66), .B(n2188), .S0(n3102), .Y(n1305) );
  MXI2XL U1340 ( .A(n67), .B(n2186), .S0(n3102), .Y(n1304) );
  MXI2XL U1341 ( .A(n68), .B(n2184), .S0(n3102), .Y(n1303) );
  MXI2XL U1342 ( .A(n69), .B(n2180), .S0(n3102), .Y(n1302) );
  MXI2XL U1343 ( .A(n71), .B(n2178), .S0(n3102), .Y(n1301) );
  MXI2XL U1344 ( .A(n72), .B(n2176), .S0(n3102), .Y(n1300) );
  MXI2XL U1345 ( .A(n73), .B(n2174), .S0(n3102), .Y(n1299) );
  MXI2XL U1346 ( .A(n74), .B(n2172), .S0(n3102), .Y(n1298) );
  MXI2XL U1347 ( .A(n75), .B(n2170), .S0(n3102), .Y(n1297) );
  MXI2XL U1348 ( .A(n76), .B(n2168), .S0(n3102), .Y(n1296) );
  MXI2XL U1349 ( .A(n77), .B(n2166), .S0(n3102), .Y(n1295) );
  MXI2XL U1350 ( .A(n78), .B(n2164), .S0(n3102), .Y(n1294) );
  MXI2XL U1351 ( .A(n79), .B(n2162), .S0(n3102), .Y(n1293) );
  MXI2XL U1352 ( .A(n80), .B(n2158), .S0(n3102), .Y(n1292) );
  MXI2XL U1353 ( .A(n81), .B(n2156), .S0(n3102), .Y(n1291) );
  MXI2XL U1354 ( .A(n82), .B(n2204), .S0(n3104), .Y(n1290) );
  MXI2XL U1355 ( .A(n83), .B(n2182), .S0(n3104), .Y(n1289) );
  MXI2XL U1356 ( .A(n84), .B(n2160), .S0(n3104), .Y(n1288) );
  MXI2XL U1357 ( .A(n85), .B(n2154), .S0(n3104), .Y(n1287) );
  MXI2XL U1358 ( .A(n86), .B(n2152), .S0(n3104), .Y(n1286) );
  MXI2XL U1359 ( .A(n87), .B(n2150), .S0(n3104), .Y(n1285) );
  MXI2XL U1360 ( .A(n88), .B(n2148), .S0(n3104), .Y(n1284) );
  MXI2XL U1361 ( .A(n89), .B(n2146), .S0(n3104), .Y(n1283) );
  MXI2XL U1362 ( .A(n90), .B(n2144), .S0(n3104), .Y(n1282) );
  MXI2XL U1363 ( .A(n91), .B(n2142), .S0(n3104), .Y(n1281) );
  MXI2XL U1364 ( .A(n92), .B(n2202), .S0(n3104), .Y(n1280) );
  MXI2XL U1365 ( .A(n93), .B(n2200), .S0(n3104), .Y(n1279) );
  MXI2XL U1366 ( .A(n94), .B(n2198), .S0(n3104), .Y(n1278) );
  MXI2XL U1367 ( .A(n95), .B(n2196), .S0(n3104), .Y(n1277) );
  MXI2XL U1368 ( .A(n96), .B(n2194), .S0(n3104), .Y(n1276) );
  MXI2XL U1369 ( .A(n97), .B(n2192), .S0(n3104), .Y(n1275) );
  MXI2XL U1370 ( .A(n98), .B(n2190), .S0(n3104), .Y(n1274) );
  MXI2XL U1371 ( .A(n99), .B(n2188), .S0(n3104), .Y(n1273) );
  MXI2XL U1372 ( .A(n100), .B(n2186), .S0(n3104), .Y(n1272) );
  MXI2XL U1373 ( .A(n101), .B(n2184), .S0(n3104), .Y(n1271) );
  MXI2XL U1374 ( .A(n102), .B(n2180), .S0(n3104), .Y(n1270) );
  MXI2XL U1375 ( .A(n103), .B(n2178), .S0(n3104), .Y(n1269) );
  MXI2XL U1376 ( .A(n104), .B(n2176), .S0(n3104), .Y(n1268) );
  MXI2XL U1377 ( .A(n105), .B(n2174), .S0(n3104), .Y(n1267) );
  MXI2XL U1378 ( .A(n106), .B(n2172), .S0(n3104), .Y(n1266) );
  MXI2XL U1379 ( .A(n107), .B(n2170), .S0(n3104), .Y(n1265) );
  MXI2XL U1380 ( .A(n108), .B(n2168), .S0(n3104), .Y(n1264) );
  MXI2XL U1381 ( .A(n109), .B(n2166), .S0(n3104), .Y(n1263) );
  MXI2XL U1382 ( .A(n110), .B(n2164), .S0(n3104), .Y(n1262) );
  MXI2XL U1383 ( .A(n111), .B(n2162), .S0(n3104), .Y(n1261) );
  MXI2XL U1384 ( .A(n112), .B(n2158), .S0(n3104), .Y(n1260) );
  MXI2XL U1385 ( .A(n113), .B(n2156), .S0(n3104), .Y(n1259) );
  MXI2XL U1386 ( .A(n114), .B(n2204), .S0(n3105), .Y(n1258) );
  MXI2XL U1387 ( .A(n115), .B(n2182), .S0(n3105), .Y(n1257) );
  MXI2XL U1388 ( .A(n116), .B(n2160), .S0(n3105), .Y(n1256) );
  MXI2XL U1389 ( .A(n117), .B(n2154), .S0(n3105), .Y(n1255) );
  MXI2XL U1390 ( .A(n118), .B(n2152), .S0(n3105), .Y(n1254) );
  MXI2XL U1391 ( .A(n119), .B(n2150), .S0(n3105), .Y(n1253) );
  MXI2XL U1392 ( .A(n120), .B(n2148), .S0(n3105), .Y(n1252) );
  MXI2XL U1393 ( .A(n121), .B(n2146), .S0(n3105), .Y(n1251) );
  MXI2XL U1394 ( .A(n122), .B(n2144), .S0(n3105), .Y(n1250) );
  MXI2XL U1395 ( .A(n123), .B(n2142), .S0(n3105), .Y(n1249) );
  MXI2XL U1396 ( .A(n124), .B(n2202), .S0(n3105), .Y(n1248) );
  MXI2XL U1397 ( .A(n125), .B(n2200), .S0(n3105), .Y(n1247) );
  MXI2XL U1398 ( .A(n126), .B(n2198), .S0(n3105), .Y(n1246) );
  MXI2XL U1399 ( .A(n127), .B(n2196), .S0(n3105), .Y(n1245) );
  MXI2XL U1400 ( .A(n128), .B(n2194), .S0(n3105), .Y(n1244) );
  MXI2XL U1401 ( .A(n129), .B(n2192), .S0(n3105), .Y(n1243) );
  MXI2XL U1402 ( .A(n130), .B(n2190), .S0(n3105), .Y(n1242) );
  MXI2XL U1403 ( .A(n131), .B(n2188), .S0(n3105), .Y(n1241) );
  MXI2XL U1404 ( .A(n132), .B(n2186), .S0(n3105), .Y(n1240) );
  MXI2XL U1405 ( .A(n133), .B(n2184), .S0(n3105), .Y(n1239) );
  MXI2XL U1406 ( .A(n134), .B(n2180), .S0(n3105), .Y(n1238) );
  MXI2XL U1407 ( .A(n135), .B(n2178), .S0(n3105), .Y(n1237) );
  MXI2XL U1408 ( .A(n136), .B(n2176), .S0(n3105), .Y(n1236) );
  MXI2XL U1409 ( .A(n137), .B(n2174), .S0(n3105), .Y(n1235) );
  MXI2XL U1410 ( .A(n138), .B(n2172), .S0(n3105), .Y(n1234) );
  MXI2XL U1411 ( .A(n139), .B(n2170), .S0(n3105), .Y(n1233) );
  MXI2XL U1412 ( .A(n140), .B(n2168), .S0(n3105), .Y(n1232) );
  MXI2XL U1413 ( .A(n141), .B(n2166), .S0(n3105), .Y(n1231) );
  MXI2XL U1414 ( .A(n142), .B(n2164), .S0(n3105), .Y(n1230) );
  MXI2XL U1415 ( .A(n143), .B(n2162), .S0(n3105), .Y(n1229) );
  MXI2XL U1416 ( .A(n144), .B(n2158), .S0(n3105), .Y(n1228) );
  MXI2XL U1417 ( .A(n145), .B(n2156), .S0(n3105), .Y(n1227) );
  MXI2XL U1418 ( .A(n146), .B(n2204), .S0(n3106), .Y(n1226) );
  MXI2XL U1419 ( .A(n147), .B(n2182), .S0(n3106), .Y(n1225) );
  MXI2XL U1420 ( .A(n148), .B(n2160), .S0(n3106), .Y(n1224) );
  MXI2XL U1421 ( .A(n149), .B(n2154), .S0(n3106), .Y(n1223) );
  MXI2XL U1422 ( .A(n150), .B(n2152), .S0(n3106), .Y(n1222) );
  MXI2XL U1423 ( .A(n151), .B(n2150), .S0(n3106), .Y(n1221) );
  MXI2XL U1424 ( .A(n152), .B(n2148), .S0(n3106), .Y(n1220) );
  MXI2XL U1425 ( .A(n153), .B(n2146), .S0(n3106), .Y(n1219) );
  MXI2XL U1426 ( .A(n154), .B(n2144), .S0(n3106), .Y(n1218) );
  MXI2XL U1427 ( .A(n155), .B(n2142), .S0(n3106), .Y(n1217) );
  MXI2XL U1428 ( .A(n156), .B(n2202), .S0(n3106), .Y(n1216) );
  MXI2XL U1429 ( .A(n157), .B(n2200), .S0(n3106), .Y(n1215) );
  MXI2XL U1430 ( .A(n158), .B(n2198), .S0(n3106), .Y(n1214) );
  MXI2XL U1431 ( .A(n159), .B(n2196), .S0(n3106), .Y(n1213) );
  MXI2XL U1432 ( .A(n160), .B(n2194), .S0(n3106), .Y(n1212) );
  MXI2XL U1433 ( .A(n161), .B(n2192), .S0(n3106), .Y(n1211) );
  MXI2XL U1434 ( .A(n162), .B(n2190), .S0(n3106), .Y(n1210) );
  MXI2XL U1435 ( .A(n163), .B(n2188), .S0(n3106), .Y(n1209) );
  MXI2XL U1436 ( .A(n164), .B(n2186), .S0(n3106), .Y(n1208) );
  MXI2XL U1437 ( .A(n165), .B(n2184), .S0(n3106), .Y(n1207) );
  MXI2XL U1438 ( .A(n166), .B(n2180), .S0(n3106), .Y(n1206) );
  MXI2XL U1439 ( .A(n167), .B(n2178), .S0(n3106), .Y(n1205) );
  MXI2XL U1440 ( .A(n168), .B(n2176), .S0(n3106), .Y(n1204) );
  MXI2XL U1441 ( .A(n169), .B(n2174), .S0(n3106), .Y(n1203) );
  MXI2XL U1442 ( .A(n170), .B(n2172), .S0(n3106), .Y(n1202) );
  MXI2XL U1443 ( .A(n171), .B(n2170), .S0(n3106), .Y(n1201) );
  MXI2XL U1444 ( .A(n172), .B(n2168), .S0(n3106), .Y(n1200) );
  MXI2XL U1445 ( .A(n173), .B(n2166), .S0(n3106), .Y(n1199) );
  MXI2XL U1446 ( .A(n174), .B(n2164), .S0(n3106), .Y(n1198) );
  MXI2XL U1447 ( .A(n175), .B(n2162), .S0(n3106), .Y(n1197) );
  MXI2XL U1448 ( .A(n176), .B(n2158), .S0(n3106), .Y(n1196) );
  MXI2XL U1449 ( .A(n177), .B(n2156), .S0(n3106), .Y(n1195) );
  MXI2XL U1450 ( .A(n178), .B(n2204), .S0(n3108), .Y(n1194) );
  MXI2XL U1451 ( .A(n179), .B(n2182), .S0(n3108), .Y(n1193) );
  MXI2XL U1452 ( .A(n180), .B(n2160), .S0(n3108), .Y(n1192) );
  MXI2XL U1453 ( .A(n181), .B(n2154), .S0(n3108), .Y(n1191) );
  MXI2XL U1454 ( .A(n182), .B(n2152), .S0(n3108), .Y(n1190) );
  MXI2XL U1455 ( .A(n183), .B(n2150), .S0(n3108), .Y(n1189) );
  MXI2XL U1456 ( .A(n184), .B(n2148), .S0(n3108), .Y(n1188) );
  MXI2XL U1457 ( .A(n185), .B(n2146), .S0(n3108), .Y(n1187) );
  MXI2XL U1458 ( .A(n186), .B(n2144), .S0(n3108), .Y(n1186) );
  MXI2XL U1459 ( .A(n187), .B(n2142), .S0(n3108), .Y(n1185) );
  MXI2XL U1460 ( .A(n188), .B(n2202), .S0(n3108), .Y(n1184) );
  MXI2XL U1461 ( .A(n189), .B(n2200), .S0(n3108), .Y(n1183) );
  MXI2XL U1462 ( .A(n190), .B(n2198), .S0(n3108), .Y(n1182) );
  MXI2XL U1463 ( .A(n191), .B(n2196), .S0(n3108), .Y(n1181) );
  MXI2XL U1464 ( .A(n192), .B(n2194), .S0(n3108), .Y(n1180) );
  MXI2XL U1465 ( .A(n193), .B(n2192), .S0(n3108), .Y(n1179) );
  MXI2XL U1466 ( .A(n194), .B(n2190), .S0(n3108), .Y(n1178) );
  MXI2XL U1467 ( .A(n195), .B(n2188), .S0(n3108), .Y(n1177) );
  MXI2XL U1468 ( .A(n196), .B(n2186), .S0(n3108), .Y(n1176) );
  MXI2XL U1469 ( .A(n197), .B(n2184), .S0(n3108), .Y(n1175) );
  MXI2XL U1470 ( .A(n198), .B(n2180), .S0(n3108), .Y(n1174) );
  MXI2XL U1471 ( .A(n199), .B(n2178), .S0(n3108), .Y(n1173) );
  MXI2XL U1472 ( .A(n200), .B(n2176), .S0(n3108), .Y(n1172) );
  MXI2XL U1473 ( .A(n201), .B(n2174), .S0(n3108), .Y(n1171) );
  MXI2XL U1474 ( .A(n202), .B(n2172), .S0(n3108), .Y(n1170) );
  MXI2XL U1475 ( .A(n203), .B(n2170), .S0(n3108), .Y(n1169) );
  MXI2XL U1476 ( .A(n204), .B(n2168), .S0(n3108), .Y(n1168) );
  MXI2XL U1477 ( .A(n205), .B(n2166), .S0(n3108), .Y(n1167) );
  MXI2XL U1478 ( .A(n206), .B(n2164), .S0(n3108), .Y(n1166) );
  MXI2XL U1479 ( .A(n207), .B(n2162), .S0(n3108), .Y(n1165) );
  MXI2XL U1480 ( .A(n208), .B(n2158), .S0(n3108), .Y(n1164) );
  MXI2XL U1481 ( .A(n209), .B(n2156), .S0(n3108), .Y(n1163) );
  MXI2XL U1482 ( .A(n210), .B(n2204), .S0(n3111), .Y(n1162) );
  MXI2XL U1483 ( .A(n211), .B(n2182), .S0(n3111), .Y(n1161) );
  MXI2XL U1484 ( .A(n212), .B(n2160), .S0(n3111), .Y(n1160) );
  MXI2XL U1485 ( .A(n213), .B(n2154), .S0(n3111), .Y(n1159) );
  MXI2XL U1486 ( .A(n214), .B(n2152), .S0(n3111), .Y(n1158) );
  MXI2XL U1487 ( .A(n215), .B(n2150), .S0(n3111), .Y(n1157) );
  MXI2XL U1488 ( .A(n216), .B(n2148), .S0(n3111), .Y(n1156) );
  MXI2XL U1489 ( .A(n217), .B(n2146), .S0(n3111), .Y(n1155) );
  MXI2XL U1490 ( .A(n218), .B(n2144), .S0(n3111), .Y(n1154) );
  MXI2XL U1491 ( .A(n219), .B(n2142), .S0(n3111), .Y(n1153) );
  MXI2XL U1492 ( .A(n220), .B(n2202), .S0(n3111), .Y(n1152) );
  MXI2XL U1493 ( .A(n221), .B(n2200), .S0(n3111), .Y(n1151) );
  MXI2XL U1494 ( .A(n222), .B(n2198), .S0(n3111), .Y(n1150) );
  MXI2XL U1495 ( .A(n223), .B(n2196), .S0(n3111), .Y(n1149) );
  MXI2XL U1496 ( .A(n224), .B(n2194), .S0(n3111), .Y(n1148) );
  MXI2XL U1497 ( .A(n225), .B(n2192), .S0(n3111), .Y(n1147) );
  MXI2XL U1498 ( .A(n226), .B(n2190), .S0(n3111), .Y(n1146) );
  MXI2XL U1499 ( .A(n227), .B(n2188), .S0(n3111), .Y(n1145) );
  MXI2XL U1500 ( .A(n228), .B(n2186), .S0(n3111), .Y(n1144) );
  MXI2XL U1501 ( .A(n229), .B(n2184), .S0(n3111), .Y(n1143) );
  MXI2XL U1502 ( .A(n230), .B(n2180), .S0(n3111), .Y(n1142) );
  MXI2XL U1503 ( .A(n231), .B(n2178), .S0(n3111), .Y(n1141) );
  MXI2XL U1504 ( .A(n232), .B(n2176), .S0(n3111), .Y(n1140) );
  MXI2XL U1505 ( .A(n233), .B(n2174), .S0(n3111), .Y(n1139) );
  MXI2XL U1506 ( .A(n234), .B(n2172), .S0(n3111), .Y(n1138) );
  MXI2XL U1507 ( .A(n235), .B(n2170), .S0(n3111), .Y(n1137) );
  MXI2XL U1508 ( .A(n236), .B(n2168), .S0(n3111), .Y(n1136) );
  MXI2XL U1509 ( .A(n237), .B(n2166), .S0(n3111), .Y(n1135) );
  MXI2XL U1510 ( .A(n238), .B(n2164), .S0(n3111), .Y(n1134) );
  MXI2XL U1511 ( .A(n239), .B(n2162), .S0(n3111), .Y(n1133) );
  MXI2XL U1512 ( .A(n240), .B(n2158), .S0(n3111), .Y(n1132) );
  MXI2XL U1513 ( .A(n241), .B(n2156), .S0(n3111), .Y(n1131) );
  MXI2XL U1514 ( .A(n242), .B(n2204), .S0(n3112), .Y(n1130) );
  MXI2XL U1515 ( .A(n243), .B(n2182), .S0(n3112), .Y(n1129) );
  MXI2XL U1516 ( .A(n244), .B(n2160), .S0(n3112), .Y(n1128) );
  MXI2XL U1517 ( .A(n245), .B(n2154), .S0(n3112), .Y(n1127) );
  MXI2XL U1518 ( .A(n246), .B(n2152), .S0(n3112), .Y(n1126) );
  MXI2XL U1519 ( .A(n247), .B(n2150), .S0(n3112), .Y(n1125) );
  MXI2XL U1520 ( .A(n248), .B(n2148), .S0(n3112), .Y(n1124) );
  MXI2XL U1521 ( .A(n249), .B(n2146), .S0(n3112), .Y(n1123) );
  MXI2XL U1522 ( .A(n250), .B(n2144), .S0(n3112), .Y(n1122) );
  MXI2XL U1523 ( .A(n251), .B(n2142), .S0(n3112), .Y(n1121) );
  MXI2XL U1524 ( .A(n252), .B(n2202), .S0(n3112), .Y(n1120) );
  MXI2XL U1525 ( .A(n253), .B(n2200), .S0(n3112), .Y(n1119) );
  MXI2XL U1526 ( .A(n254), .B(n2198), .S0(n3112), .Y(n1118) );
  MXI2XL U1527 ( .A(n255), .B(n2196), .S0(n3112), .Y(n1117) );
  MXI2XL U1528 ( .A(n256), .B(n2194), .S0(n3112), .Y(n1116) );
  MXI2XL U1529 ( .A(n257), .B(n2192), .S0(n3112), .Y(n1115) );
  MXI2XL U1530 ( .A(n258), .B(n2190), .S0(n3112), .Y(n1114) );
  MXI2XL U1531 ( .A(n259), .B(n2188), .S0(n3112), .Y(n1113) );
  MXI2XL U1532 ( .A(n260), .B(n2186), .S0(n3112), .Y(n1112) );
  MXI2XL U1533 ( .A(n261), .B(n2184), .S0(n3112), .Y(n1111) );
  MXI2XL U1534 ( .A(n262), .B(n2180), .S0(n3112), .Y(n1110) );
  MXI2XL U1535 ( .A(n263), .B(n2178), .S0(n3112), .Y(n1109) );
  MXI2XL U1536 ( .A(n264), .B(n2176), .S0(n3112), .Y(n1108) );
  MXI2XL U1537 ( .A(n265), .B(n2174), .S0(n3112), .Y(n1107) );
  MXI2XL U1538 ( .A(n266), .B(n2172), .S0(n3112), .Y(n1106) );
  MXI2XL U1539 ( .A(n267), .B(n2170), .S0(n3112), .Y(n1105) );
  MXI2XL U1540 ( .A(n268), .B(n2168), .S0(n3112), .Y(n1104) );
  MXI2XL U1541 ( .A(n269), .B(n2166), .S0(n3112), .Y(n1103) );
  MXI2XL U1542 ( .A(n270), .B(n2164), .S0(n3112), .Y(n1102) );
  MXI2XL U1543 ( .A(n271), .B(n2162), .S0(n3112), .Y(n1101) );
  MXI2XL U1544 ( .A(n272), .B(n2158), .S0(n3112), .Y(n1100) );
  MXI2XL U1545 ( .A(n273), .B(n2156), .S0(n3112), .Y(n1099) );
  MXI2XL U1546 ( .A(n274), .B(n2204), .S0(n3113), .Y(n1098) );
  MXI2XL U1547 ( .A(n275), .B(n2182), .S0(n3113), .Y(n1097) );
  MXI2XL U1548 ( .A(n276), .B(n2160), .S0(n3113), .Y(n1096) );
  MXI2XL U1549 ( .A(n277), .B(n2154), .S0(n3113), .Y(n1095) );
  MXI2XL U1550 ( .A(n278), .B(n2152), .S0(n3113), .Y(n1094) );
  MXI2XL U1551 ( .A(n279), .B(n2150), .S0(n3113), .Y(n1093) );
  MXI2XL U1552 ( .A(n280), .B(n2148), .S0(n3113), .Y(n1092) );
  MXI2XL U1553 ( .A(n281), .B(n2146), .S0(n3113), .Y(n1091) );
  MXI2XL U1554 ( .A(n282), .B(n2144), .S0(n3113), .Y(n1090) );
  MXI2XL U1555 ( .A(n283), .B(n2142), .S0(n3113), .Y(n1089) );
  MXI2XL U1556 ( .A(n284), .B(n2202), .S0(n3113), .Y(n1088) );
  MXI2XL U1557 ( .A(n285), .B(n2200), .S0(n3113), .Y(n1087) );
  MXI2XL U1558 ( .A(n286), .B(n2198), .S0(n3113), .Y(n1086) );
  MXI2XL U1559 ( .A(n287), .B(n2196), .S0(n3113), .Y(n1085) );
  MXI2XL U1560 ( .A(n288), .B(n2194), .S0(n3113), .Y(n1084) );
  MXI2XL U1561 ( .A(n289), .B(n2192), .S0(n3113), .Y(n1083) );
  MXI2XL U1562 ( .A(n290), .B(n2190), .S0(n3113), .Y(n1082) );
  MXI2XL U1563 ( .A(n291), .B(n2188), .S0(n3113), .Y(n1081) );
  MXI2XL U1564 ( .A(n292), .B(n2186), .S0(n3113), .Y(n1080) );
  MXI2XL U1565 ( .A(n293), .B(n2184), .S0(n3113), .Y(n1079) );
  MXI2XL U1566 ( .A(n294), .B(n2180), .S0(n3113), .Y(n1078) );
  MXI2XL U1567 ( .A(n295), .B(n2178), .S0(n3113), .Y(n1077) );
  MXI2XL U1568 ( .A(n296), .B(n2176), .S0(n3113), .Y(n1076) );
  MXI2XL U1569 ( .A(n297), .B(n2174), .S0(n3113), .Y(n1075) );
  MXI2XL U1570 ( .A(n298), .B(n2172), .S0(n3113), .Y(n1074) );
  MXI2XL U1571 ( .A(n1355), .B(n2170), .S0(n3113), .Y(n1073) );
  MXI2XL U1572 ( .A(n1356), .B(n2168), .S0(n3113), .Y(n1072) );
  MXI2XL U1573 ( .A(n1357), .B(n2166), .S0(n3113), .Y(n1071) );
  MXI2XL U1574 ( .A(n1358), .B(n2164), .S0(n3113), .Y(n1070) );
  MXI2XL U1575 ( .A(n1359), .B(n2162), .S0(n3113), .Y(n1069) );
  MXI2XL U1576 ( .A(n1360), .B(n2158), .S0(n3113), .Y(n1068) );
  MXI2XL U1577 ( .A(n1361), .B(n2156), .S0(n3113), .Y(n1067) );
  MXI2XL U1578 ( .A(n1362), .B(n2204), .S0(n3114), .Y(n1066) );
  MXI2XL U1579 ( .A(n1363), .B(n2182), .S0(n3114), .Y(n1065) );
  MXI2XL U1580 ( .A(n1364), .B(n2160), .S0(n3114), .Y(n1064) );
  MXI2XL U1581 ( .A(n1365), .B(n2154), .S0(n3114), .Y(n1063) );
  MXI2XL U1582 ( .A(n1366), .B(n2152), .S0(n3114), .Y(n1062) );
  MXI2XL U1583 ( .A(n1367), .B(n2150), .S0(n3114), .Y(n1061) );
  MXI2XL U1584 ( .A(n1368), .B(n2148), .S0(n3114), .Y(n1060) );
  MXI2XL U1585 ( .A(n1369), .B(n2146), .S0(n3114), .Y(n1059) );
  MXI2XL U1586 ( .A(n1370), .B(n2144), .S0(n3114), .Y(n1058) );
  MXI2XL U1587 ( .A(n1371), .B(n2142), .S0(n3114), .Y(n1057) );
  MXI2XL U1588 ( .A(n1372), .B(n2202), .S0(n3114), .Y(n1056) );
  MXI2XL U1589 ( .A(n1373), .B(n2200), .S0(n3114), .Y(n1055) );
  MXI2XL U1590 ( .A(n1374), .B(n2198), .S0(n3114), .Y(n1054) );
  MXI2XL U1591 ( .A(n1375), .B(n2196), .S0(n3114), .Y(n1053) );
  MXI2XL U1592 ( .A(n1376), .B(n2194), .S0(n3114), .Y(n1052) );
  MXI2XL U1593 ( .A(n1377), .B(n2192), .S0(n3114), .Y(n1051) );
  MXI2XL U1594 ( .A(n1378), .B(n2190), .S0(n3114), .Y(n1050) );
  MXI2XL U1595 ( .A(n1379), .B(n2188), .S0(n3114), .Y(n1049) );
  MXI2XL U1596 ( .A(n1380), .B(n2186), .S0(n3114), .Y(n1048) );
  MXI2XL U1597 ( .A(n1381), .B(n2184), .S0(n3114), .Y(n1047) );
  MXI2XL U1598 ( .A(n1382), .B(n2180), .S0(n3114), .Y(n1046) );
  MXI2XL U1599 ( .A(n1383), .B(n2178), .S0(n3114), .Y(n1045) );
  MXI2XL U1600 ( .A(n1384), .B(n2176), .S0(n3114), .Y(n1044) );
  MXI2XL U1601 ( .A(n1385), .B(n2174), .S0(n3114), .Y(n1043) );
  MXI2XL U1602 ( .A(n1386), .B(n2172), .S0(n3114), .Y(n1042) );
  MXI2XL U1603 ( .A(n1387), .B(n2170), .S0(n3114), .Y(n1041) );
  MXI2XL U1604 ( .A(n1388), .B(n2168), .S0(n3114), .Y(n1040) );
  MXI2XL U1605 ( .A(n1389), .B(n2166), .S0(n3114), .Y(n1039) );
  MXI2XL U1606 ( .A(n1390), .B(n2164), .S0(n3114), .Y(n1038) );
  MXI2XL U1607 ( .A(n1391), .B(n2162), .S0(n3114), .Y(n1037) );
  MXI2XL U1608 ( .A(n1392), .B(n2158), .S0(n3114), .Y(n1036) );
  MXI2XL U1609 ( .A(n1393), .B(n2156), .S0(n3114), .Y(n1035) );
  MXI2XL U1610 ( .A(n1394), .B(n2204), .S0(n3115), .Y(n1034) );
  MXI2XL U1611 ( .A(n1395), .B(n2182), .S0(n3115), .Y(n1033) );
  MXI2XL U1612 ( .A(n1396), .B(n2160), .S0(n3115), .Y(n1032) );
  MXI2XL U1613 ( .A(n1397), .B(n2154), .S0(n3115), .Y(n1031) );
  MXI2XL U1614 ( .A(n1398), .B(n2152), .S0(n3115), .Y(n1030) );
  MXI2XL U1615 ( .A(n1399), .B(n2150), .S0(n3115), .Y(n1029) );
  MXI2XL U1616 ( .A(n1400), .B(n2148), .S0(n3115), .Y(n1028) );
  MXI2XL U1617 ( .A(n1401), .B(n2146), .S0(n3115), .Y(n1027) );
  MXI2XL U1618 ( .A(n1402), .B(n2144), .S0(n3115), .Y(n1026) );
  MXI2XL U1619 ( .A(n1403), .B(n2142), .S0(n3115), .Y(n1025) );
  MXI2XL U1620 ( .A(n1404), .B(n2202), .S0(n3115), .Y(n1024) );
  MXI2XL U1621 ( .A(n1405), .B(n2200), .S0(n3115), .Y(n1023) );
  MXI2XL U1622 ( .A(n1406), .B(n2198), .S0(n3115), .Y(n1022) );
  MXI2XL U1623 ( .A(n1407), .B(n2196), .S0(n3115), .Y(n1021) );
  MXI2XL U1624 ( .A(n1408), .B(n2194), .S0(n3115), .Y(n1020) );
  MXI2XL U1625 ( .A(n1409), .B(n2192), .S0(n3115), .Y(n1019) );
  MXI2XL U1626 ( .A(n1410), .B(n2190), .S0(n3115), .Y(n1018) );
  MXI2XL U1627 ( .A(n1411), .B(n2188), .S0(n3115), .Y(n1017) );
  MXI2XL U1628 ( .A(n1412), .B(n2186), .S0(n3115), .Y(n1016) );
  MXI2XL U1629 ( .A(n1413), .B(n2184), .S0(n3115), .Y(n1015) );
  MXI2XL U1630 ( .A(n1414), .B(n2180), .S0(n3115), .Y(n1014) );
  MXI2XL U1631 ( .A(n1415), .B(n2178), .S0(n3115), .Y(n1013) );
  MXI2XL U1632 ( .A(n1416), .B(n2176), .S0(n3115), .Y(n1012) );
  MXI2XL U1633 ( .A(n1417), .B(n2174), .S0(n3115), .Y(n1011) );
  MXI2XL U1634 ( .A(n1418), .B(n2172), .S0(n3115), .Y(n1010) );
  MXI2XL U1635 ( .A(n1419), .B(n2170), .S0(n3115), .Y(n1009) );
  MXI2XL U1636 ( .A(n1420), .B(n2168), .S0(n3115), .Y(n1008) );
  MXI2XL U1637 ( .A(n1421), .B(n2166), .S0(n3115), .Y(n1007) );
  MXI2XL U1638 ( .A(n1422), .B(n2164), .S0(n3115), .Y(n1006) );
  MXI2XL U1639 ( .A(n1423), .B(n2162), .S0(n3115), .Y(n1005) );
  MXI2XL U1640 ( .A(n1424), .B(n2158), .S0(n3115), .Y(n1004) );
  MXI2XL U1641 ( .A(n1425), .B(n2156), .S0(n3115), .Y(n1003) );
  MXI2XL U1642 ( .A(n1426), .B(n2204), .S0(n2991), .Y(n1002) );
  MXI2XL U1643 ( .A(n1427), .B(n2182), .S0(n2991), .Y(n1001) );
  MXI2XL U1644 ( .A(n1428), .B(n2160), .S0(n2991), .Y(n1000) );
  MXI2XL U1645 ( .A(n1429), .B(n2154), .S0(n2991), .Y(n999) );
  MXI2XL U1646 ( .A(n1430), .B(n2152), .S0(n2991), .Y(n998) );
  MXI2XL U1647 ( .A(n1431), .B(n2150), .S0(n2991), .Y(n997) );
  MXI2XL U1648 ( .A(n1432), .B(n2148), .S0(n2991), .Y(n996) );
  MXI2XL U1649 ( .A(n1433), .B(n2146), .S0(n2991), .Y(n995) );
  MXI2XL U1650 ( .A(n1434), .B(n2144), .S0(n2991), .Y(n994) );
  MXI2XL U1651 ( .A(n1435), .B(n2142), .S0(n2991), .Y(n993) );
  MXI2XL U1652 ( .A(n1436), .B(n2202), .S0(n2991), .Y(n992) );
  MXI2XL U1653 ( .A(n1437), .B(n2200), .S0(n2991), .Y(n991) );
  MXI2XL U1654 ( .A(n1438), .B(n2198), .S0(n2991), .Y(n990) );
  MXI2XL U1655 ( .A(n1439), .B(n2196), .S0(n2991), .Y(n989) );
  MXI2XL U1656 ( .A(n1440), .B(n2194), .S0(n2991), .Y(n988) );
  MXI2XL U1657 ( .A(n1441), .B(n2192), .S0(n2991), .Y(n987) );
  MXI2XL U1658 ( .A(n1442), .B(n2190), .S0(n2991), .Y(n986) );
  MXI2XL U1659 ( .A(n1443), .B(n2188), .S0(n2991), .Y(n985) );
  MXI2XL U1660 ( .A(n1444), .B(n2186), .S0(n2991), .Y(n984) );
  MXI2XL U1661 ( .A(n1445), .B(n2184), .S0(n2991), .Y(n983) );
  MXI2XL U1662 ( .A(n1446), .B(n2180), .S0(n2991), .Y(n982) );
  MXI2XL U1663 ( .A(n1447), .B(n2178), .S0(n2991), .Y(n981) );
  MXI2XL U1664 ( .A(n1448), .B(n2176), .S0(n2991), .Y(n980) );
  MXI2XL U1665 ( .A(n1449), .B(n2174), .S0(n2991), .Y(n979) );
  MXI2XL U1666 ( .A(n1450), .B(n2172), .S0(n2991), .Y(n978) );
  MXI2XL U1667 ( .A(n1451), .B(n2170), .S0(n2991), .Y(n977) );
  MXI2XL U1668 ( .A(n1452), .B(n2168), .S0(n2991), .Y(n976) );
  MXI2XL U1669 ( .A(n1453), .B(n2166), .S0(n2991), .Y(n975) );
  MXI2XL U1670 ( .A(n1454), .B(n2164), .S0(n2991), .Y(n974) );
  MXI2XL U1671 ( .A(n1455), .B(n2162), .S0(n2991), .Y(n973) );
  MXI2XL U1672 ( .A(n1456), .B(n2158), .S0(n2991), .Y(n972) );
  MXI2XL U1673 ( .A(n1457), .B(n2156), .S0(n2991), .Y(n971) );
  MXI2XL U1674 ( .A(n1458), .B(n2204), .S0(n2992), .Y(n970) );
  MXI2XL U1675 ( .A(n1459), .B(n2182), .S0(n2992), .Y(n969) );
  MXI2XL U1676 ( .A(n1460), .B(n2160), .S0(n2992), .Y(n968) );
  MXI2XL U1677 ( .A(n1461), .B(n2154), .S0(n2992), .Y(n967) );
  MXI2XL U1678 ( .A(n1462), .B(n2152), .S0(n2992), .Y(n966) );
  MXI2XL U1679 ( .A(n1463), .B(n2150), .S0(n2992), .Y(n965) );
  MXI2XL U1680 ( .A(n1464), .B(n2148), .S0(n2992), .Y(n964) );
  MXI2XL U1681 ( .A(n1465), .B(n2146), .S0(n2992), .Y(n963) );
  MXI2XL U1682 ( .A(n1466), .B(n2144), .S0(n2992), .Y(n962) );
  MXI2XL U1683 ( .A(n1467), .B(n2142), .S0(n2992), .Y(n961) );
  MXI2XL U1684 ( .A(n1468), .B(n2202), .S0(n2992), .Y(n960) );
  MXI2XL U1685 ( .A(n1469), .B(n2200), .S0(n2992), .Y(n959) );
  MXI2XL U1686 ( .A(n1470), .B(n2198), .S0(n2992), .Y(n958) );
  MXI2XL U1687 ( .A(n1471), .B(n2196), .S0(n2992), .Y(n957) );
  MXI2XL U1688 ( .A(n1472), .B(n2194), .S0(n2992), .Y(n956) );
  MXI2XL U1689 ( .A(n1473), .B(n2192), .S0(n2992), .Y(n955) );
  MXI2XL U1690 ( .A(n1474), .B(n2190), .S0(n2992), .Y(n954) );
  MXI2XL U1691 ( .A(n1475), .B(n2188), .S0(n2992), .Y(n953) );
  MXI2XL U1692 ( .A(n1476), .B(n2186), .S0(n2992), .Y(n952) );
  MXI2XL U1693 ( .A(n1477), .B(n2184), .S0(n2992), .Y(n951) );
  MXI2XL U1694 ( .A(n1478), .B(n2180), .S0(n2992), .Y(n950) );
  MXI2XL U1695 ( .A(n1479), .B(n2178), .S0(n2992), .Y(n949) );
  MXI2XL U1696 ( .A(n1480), .B(n2176), .S0(n2992), .Y(n948) );
  MXI2XL U1697 ( .A(n1481), .B(n2174), .S0(n2992), .Y(n947) );
  MXI2XL U1698 ( .A(n1482), .B(n2172), .S0(n2992), .Y(n946) );
  MXI2XL U1699 ( .A(n1483), .B(n2170), .S0(n2992), .Y(n945) );
  MXI2XL U1700 ( .A(n1484), .B(n2168), .S0(n2992), .Y(n944) );
  MXI2XL U1701 ( .A(n1485), .B(n2166), .S0(n2992), .Y(n943) );
  MXI2XL U1702 ( .A(n1486), .B(n2164), .S0(n2992), .Y(n942) );
  MXI2XL U1703 ( .A(n1487), .B(n2162), .S0(n2992), .Y(n941) );
  MXI2XL U1704 ( .A(n1488), .B(n2158), .S0(n2992), .Y(n940) );
  MXI2XL U1705 ( .A(n1489), .B(n2156), .S0(n2992), .Y(n939) );
  MXI2XL U1706 ( .A(n1490), .B(n2204), .S0(n2995), .Y(n938) );
  MXI2XL U1707 ( .A(n1491), .B(n2182), .S0(n2995), .Y(n937) );
  MXI2XL U1708 ( .A(n1492), .B(n2160), .S0(n2995), .Y(n936) );
  MXI2XL U1709 ( .A(n1493), .B(n2154), .S0(n2995), .Y(n935) );
  MXI2XL U1710 ( .A(n1494), .B(n2152), .S0(n2995), .Y(n934) );
  MXI2XL U1711 ( .A(n1495), .B(n2150), .S0(n2995), .Y(n933) );
  MXI2XL U1712 ( .A(n1496), .B(n2148), .S0(n2995), .Y(n932) );
  MXI2XL U1713 ( .A(n1497), .B(n2146), .S0(n2995), .Y(n931) );
  MXI2XL U1714 ( .A(n1498), .B(n2144), .S0(n2995), .Y(n930) );
  MXI2XL U1715 ( .A(n1499), .B(n2142), .S0(n2995), .Y(n929) );
  MXI2XL U1716 ( .A(n1500), .B(n2202), .S0(n2995), .Y(n928) );
  MXI2XL U1717 ( .A(n1501), .B(n2200), .S0(n2995), .Y(n927) );
  MXI2XL U1718 ( .A(n1502), .B(n2198), .S0(n2995), .Y(n926) );
  MXI2XL U1719 ( .A(n1503), .B(n2196), .S0(n2995), .Y(n925) );
  MXI2XL U1720 ( .A(n1504), .B(n2194), .S0(n2995), .Y(n924) );
  MXI2XL U1721 ( .A(n1505), .B(n2192), .S0(n2995), .Y(n923) );
  MXI2XL U1722 ( .A(n1506), .B(n2190), .S0(n2995), .Y(n922) );
  MXI2XL U1723 ( .A(n1507), .B(n2188), .S0(n2995), .Y(n921) );
  MXI2XL U1724 ( .A(n1508), .B(n2186), .S0(n2995), .Y(n920) );
  MXI2XL U1725 ( .A(n1509), .B(n2184), .S0(n2995), .Y(n919) );
  MXI2XL U1726 ( .A(n1510), .B(n2180), .S0(n2995), .Y(n918) );
  MXI2XL U1727 ( .A(n1511), .B(n2178), .S0(n2995), .Y(n917) );
  MXI2XL U1728 ( .A(n1512), .B(n2176), .S0(n2995), .Y(n916) );
  MXI2XL U1729 ( .A(n1513), .B(n2174), .S0(n2995), .Y(n915) );
  MXI2XL U1730 ( .A(n1514), .B(n2172), .S0(n2995), .Y(n914) );
  MXI2XL U1731 ( .A(n1515), .B(n2170), .S0(n2995), .Y(n913) );
  MXI2XL U1732 ( .A(n1516), .B(n2168), .S0(n2995), .Y(n912) );
  MXI2XL U1733 ( .A(n1517), .B(n2166), .S0(n2995), .Y(n911) );
  MXI2XL U1734 ( .A(n1518), .B(n2164), .S0(n2995), .Y(n910) );
  MXI2XL U1735 ( .A(n1519), .B(n2162), .S0(n2995), .Y(n909) );
  MXI2XL U1736 ( .A(n1520), .B(n2158), .S0(n2995), .Y(n908) );
  MXI2XL U1737 ( .A(n1521), .B(n2156), .S0(n2995), .Y(n907) );
  MXI2XL U1738 ( .A(n1522), .B(n2204), .S0(n2997), .Y(n906) );
  MXI2XL U1739 ( .A(n1523), .B(n2182), .S0(n2997), .Y(n905) );
  MXI2XL U1740 ( .A(n1524), .B(n2160), .S0(n2997), .Y(n904) );
  MXI2XL U1741 ( .A(n1525), .B(n2154), .S0(n2997), .Y(n903) );
  MXI2XL U1742 ( .A(n1526), .B(n2152), .S0(n2997), .Y(n902) );
  MXI2XL U1743 ( .A(n1527), .B(n2150), .S0(n2997), .Y(n901) );
  MXI2XL U1744 ( .A(n1528), .B(n2148), .S0(n2997), .Y(n900) );
  MXI2XL U1745 ( .A(n1529), .B(n2146), .S0(n2997), .Y(n899) );
  MXI2XL U1746 ( .A(n1530), .B(n2144), .S0(n2997), .Y(n898) );
  MXI2XL U1747 ( .A(n1531), .B(n2142), .S0(n2997), .Y(n897) );
  MXI2XL U1748 ( .A(n1532), .B(n2202), .S0(n2997), .Y(n896) );
  MXI2XL U1749 ( .A(n1533), .B(n2200), .S0(n2997), .Y(n895) );
  MXI2XL U1750 ( .A(n1534), .B(n2198), .S0(n2997), .Y(n894) );
  MXI2XL U1751 ( .A(n1535), .B(n2196), .S0(n2997), .Y(n893) );
  MXI2XL U1752 ( .A(n1536), .B(n2194), .S0(n2997), .Y(n892) );
  MXI2XL U1753 ( .A(n1537), .B(n2192), .S0(n2997), .Y(n891) );
  MXI2XL U1754 ( .A(n1538), .B(n2190), .S0(n2997), .Y(n890) );
  MXI2XL U1755 ( .A(n1539), .B(n2188), .S0(n2997), .Y(n889) );
  MXI2XL U1756 ( .A(n1540), .B(n2186), .S0(n2997), .Y(n888) );
  MXI2XL U1757 ( .A(n1541), .B(n2184), .S0(n2997), .Y(n887) );
  MXI2XL U1758 ( .A(n1542), .B(n2180), .S0(n2997), .Y(n886) );
  MXI2XL U1759 ( .A(n1543), .B(n2178), .S0(n2997), .Y(n885) );
  MXI2XL U1760 ( .A(n1544), .B(n2176), .S0(n2997), .Y(n884) );
  MXI2XL U1761 ( .A(n1545), .B(n2174), .S0(n2997), .Y(n883) );
  MXI2XL U1762 ( .A(n1546), .B(n2172), .S0(n2997), .Y(n882) );
  MXI2XL U1763 ( .A(n1547), .B(n2170), .S0(n2997), .Y(n881) );
  MXI2XL U1764 ( .A(n1548), .B(n2168), .S0(n2997), .Y(n880) );
  MXI2XL U1765 ( .A(n1549), .B(n2166), .S0(n2997), .Y(n879) );
  MXI2XL U1766 ( .A(n1550), .B(n2164), .S0(n2997), .Y(n878) );
  MXI2XL U1767 ( .A(n1551), .B(n2162), .S0(n2997), .Y(n877) );
  MXI2XL U1768 ( .A(n1552), .B(n2158), .S0(n2997), .Y(n876) );
  MXI2XL U1769 ( .A(n1553), .B(n2156), .S0(n2997), .Y(n875) );
  MXI2XL U1770 ( .A(n1554), .B(n2204), .S0(n2999), .Y(n874) );
  MXI2XL U1771 ( .A(n1555), .B(n2182), .S0(n2999), .Y(n873) );
  MXI2XL U1772 ( .A(n1556), .B(n2160), .S0(n2999), .Y(n872) );
  MXI2XL U1773 ( .A(n1557), .B(n2154), .S0(n2999), .Y(n871) );
  MXI2XL U1774 ( .A(n1558), .B(n2152), .S0(n2999), .Y(n870) );
  MXI2XL U1775 ( .A(n1559), .B(n2150), .S0(n2999), .Y(n869) );
  MXI2XL U1776 ( .A(n1560), .B(n2148), .S0(n2999), .Y(n868) );
  MXI2XL U1777 ( .A(n1561), .B(n2146), .S0(n2999), .Y(n867) );
  MXI2XL U1778 ( .A(n1562), .B(n2144), .S0(n2999), .Y(n866) );
  MXI2XL U1779 ( .A(n1563), .B(n2142), .S0(n2999), .Y(n865) );
  MXI2XL U1780 ( .A(n1564), .B(n2202), .S0(n2999), .Y(n864) );
  MXI2XL U1781 ( .A(n1565), .B(n2200), .S0(n2999), .Y(n863) );
  MXI2XL U1782 ( .A(n1566), .B(n2198), .S0(n2999), .Y(n862) );
  MXI2XL U1783 ( .A(n1567), .B(n2196), .S0(n2999), .Y(n861) );
  MXI2XL U1784 ( .A(n1568), .B(n2194), .S0(n2999), .Y(n860) );
  MXI2XL U1785 ( .A(n1569), .B(n2192), .S0(n2999), .Y(n859) );
  MXI2XL U1786 ( .A(n1570), .B(n2190), .S0(n2999), .Y(n858) );
  MXI2XL U1787 ( .A(n1571), .B(n2188), .S0(n2999), .Y(n857) );
  MXI2XL U1788 ( .A(n1572), .B(n2186), .S0(n2999), .Y(n856) );
  MXI2XL U1789 ( .A(n1573), .B(n2184), .S0(n2999), .Y(n855) );
  MXI2XL U1790 ( .A(n1574), .B(n2180), .S0(n2999), .Y(n854) );
  MXI2XL U1791 ( .A(n1575), .B(n2178), .S0(n2999), .Y(n853) );
  MXI2XL U1792 ( .A(n1576), .B(n2176), .S0(n2999), .Y(n852) );
  MXI2XL U1793 ( .A(n1577), .B(n2174), .S0(n2999), .Y(n851) );
  MXI2XL U1794 ( .A(n1578), .B(n2172), .S0(n2999), .Y(n850) );
  MXI2XL U1795 ( .A(n1579), .B(n2170), .S0(n2999), .Y(n849) );
  MXI2XL U1796 ( .A(n1580), .B(n2168), .S0(n2999), .Y(n848) );
  MXI2XL U1797 ( .A(n1581), .B(n2166), .S0(n2999), .Y(n847) );
  MXI2XL U1798 ( .A(n1582), .B(n2164), .S0(n2999), .Y(n846) );
  MXI2XL U1799 ( .A(n1583), .B(n2162), .S0(n2999), .Y(n845) );
  MXI2XL U1800 ( .A(n1584), .B(n2158), .S0(n2999), .Y(n844) );
  MXI2XL U1801 ( .A(n1585), .B(n2156), .S0(n2999), .Y(n843) );
  MXI2XL U1802 ( .A(n1586), .B(n2204), .S0(n3001), .Y(n842) );
  MXI2XL U1803 ( .A(n1587), .B(n2182), .S0(n3001), .Y(n841) );
  MXI2XL U1804 ( .A(n1588), .B(n2160), .S0(n3001), .Y(n840) );
  MXI2XL U1805 ( .A(n1589), .B(n2154), .S0(n3001), .Y(n839) );
  MXI2XL U1806 ( .A(n1590), .B(n2152), .S0(n3001), .Y(n838) );
  MXI2XL U1807 ( .A(n1591), .B(n2150), .S0(n3001), .Y(n837) );
  MXI2XL U1808 ( .A(n1592), .B(n2148), .S0(n3001), .Y(n836) );
  MXI2XL U1809 ( .A(n1593), .B(n2146), .S0(n3001), .Y(n835) );
  MXI2XL U1810 ( .A(n1594), .B(n2144), .S0(n3001), .Y(n834) );
  MXI2XL U1811 ( .A(n1595), .B(n2142), .S0(n3001), .Y(n833) );
  MXI2XL U1812 ( .A(n1596), .B(n2202), .S0(n3001), .Y(n832) );
  MXI2XL U1813 ( .A(n1597), .B(n2200), .S0(n3001), .Y(n831) );
  MXI2XL U1814 ( .A(n1598), .B(n2198), .S0(n3001), .Y(n830) );
  MXI2XL U1815 ( .A(n1599), .B(n2196), .S0(n3001), .Y(n829) );
  MXI2XL U1816 ( .A(n1600), .B(n2194), .S0(n3001), .Y(n828) );
  MXI2XL U1817 ( .A(n1601), .B(n2192), .S0(n3001), .Y(n827) );
  MXI2XL U1818 ( .A(n1602), .B(n2190), .S0(n3001), .Y(n826) );
  MXI2XL U1819 ( .A(n1603), .B(n2188), .S0(n3001), .Y(n825) );
  MXI2XL U1820 ( .A(n1604), .B(n2186), .S0(n3001), .Y(n824) );
  MXI2XL U1821 ( .A(n1605), .B(n2184), .S0(n3001), .Y(n823) );
  MXI2XL U1822 ( .A(n1606), .B(n2180), .S0(n3001), .Y(n822) );
  MXI2XL U1823 ( .A(n1607), .B(n2178), .S0(n3001), .Y(n821) );
  MXI2XL U1824 ( .A(n1608), .B(n2176), .S0(n3001), .Y(n820) );
  MXI2XL U1825 ( .A(n1609), .B(n2174), .S0(n3001), .Y(n819) );
  MXI2XL U1826 ( .A(n1610), .B(n2172), .S0(n3001), .Y(n818) );
  MXI2XL U1827 ( .A(n1611), .B(n2170), .S0(n3001), .Y(n817) );
  MXI2XL U1828 ( .A(n1612), .B(n2168), .S0(n3001), .Y(n816) );
  MXI2XL U1829 ( .A(n1613), .B(n2166), .S0(n3001), .Y(n815) );
  MXI2XL U1830 ( .A(n1614), .B(n2164), .S0(n3001), .Y(n814) );
  MXI2XL U1831 ( .A(n1615), .B(n2162), .S0(n3001), .Y(n813) );
  MXI2XL U1832 ( .A(n1616), .B(n2158), .S0(n3001), .Y(n812) );
  MXI2XL U1833 ( .A(n1617), .B(n2156), .S0(n3001), .Y(n811) );
  MXI2XL U1834 ( .A(n1618), .B(n2204), .S0(n3003), .Y(n810) );
  MXI2XL U1835 ( .A(n1619), .B(n2182), .S0(n3003), .Y(n809) );
  MXI2XL U1836 ( .A(n1620), .B(n2160), .S0(n3003), .Y(n808) );
  MXI2XL U1837 ( .A(n1621), .B(n2154), .S0(n3003), .Y(n807) );
  MXI2XL U1838 ( .A(n1622), .B(n2152), .S0(n3003), .Y(n806) );
  MXI2XL U1839 ( .A(n1623), .B(n2150), .S0(n3003), .Y(n805) );
  MXI2XL U1840 ( .A(n1624), .B(n2148), .S0(n3003), .Y(n804) );
  MXI2XL U1841 ( .A(n1625), .B(n2146), .S0(n3003), .Y(n803) );
  MXI2XL U1842 ( .A(n1626), .B(n2144), .S0(n3003), .Y(n802) );
  MXI2XL U1843 ( .A(n1627), .B(n2142), .S0(n3003), .Y(n801) );
  MXI2XL U1844 ( .A(n1628), .B(n2202), .S0(n3003), .Y(n800) );
  MXI2XL U1845 ( .A(n1629), .B(n2200), .S0(n3003), .Y(n799) );
  MXI2XL U1846 ( .A(n1630), .B(n2198), .S0(n3003), .Y(n798) );
  MXI2XL U1847 ( .A(n1631), .B(n2196), .S0(n3003), .Y(n797) );
  MXI2XL U1848 ( .A(n1632), .B(n2194), .S0(n3003), .Y(n796) );
  MXI2XL U1849 ( .A(n1633), .B(n2192), .S0(n3003), .Y(n795) );
  MXI2XL U1850 ( .A(n1634), .B(n2190), .S0(n3003), .Y(n794) );
  MXI2XL U1851 ( .A(n1635), .B(n2188), .S0(n3003), .Y(n793) );
  MXI2XL U1852 ( .A(n1636), .B(n2186), .S0(n3003), .Y(n792) );
  MXI2XL U1853 ( .A(n1637), .B(n2184), .S0(n3003), .Y(n791) );
  MXI2XL U1854 ( .A(n1638), .B(n2180), .S0(n3003), .Y(n790) );
  MXI2XL U1855 ( .A(n1639), .B(n2178), .S0(n3003), .Y(n789) );
  MXI2XL U1856 ( .A(n1640), .B(n2176), .S0(n3003), .Y(n788) );
  MXI2XL U1857 ( .A(n1641), .B(n2174), .S0(n3003), .Y(n787) );
  MXI2XL U1858 ( .A(n1642), .B(n2172), .S0(n3003), .Y(n786) );
  MXI2XL U1859 ( .A(n1643), .B(n2170), .S0(n3003), .Y(n785) );
  MXI2XL U1860 ( .A(n1644), .B(n2168), .S0(n3003), .Y(n784) );
  MXI2XL U1861 ( .A(n1645), .B(n2166), .S0(n3003), .Y(n783) );
  MXI2XL U1862 ( .A(n1646), .B(n2164), .S0(n3003), .Y(n782) );
  MXI2XL U1863 ( .A(n1647), .B(n2162), .S0(n3003), .Y(n781) );
  MXI2XL U1864 ( .A(n1648), .B(n2158), .S0(n3003), .Y(n780) );
  MXI2XL U1865 ( .A(n1649), .B(n2156), .S0(n3003), .Y(n779) );
  MXI2XL U1866 ( .A(n1650), .B(n2204), .S0(n3006), .Y(n778) );
  MXI2XL U1867 ( .A(n1651), .B(n2182), .S0(n3006), .Y(n777) );
  MXI2XL U1868 ( .A(n1652), .B(n2160), .S0(n3006), .Y(n776) );
  MXI2XL U1869 ( .A(n1653), .B(n2154), .S0(n3006), .Y(n775) );
  MXI2XL U1870 ( .A(n1654), .B(n2152), .S0(n3006), .Y(n774) );
  MXI2XL U1871 ( .A(n1655), .B(n2150), .S0(n3006), .Y(n773) );
  MXI2XL U1872 ( .A(n1656), .B(n2148), .S0(n3006), .Y(n772) );
  MXI2XL U1873 ( .A(n1657), .B(n2146), .S0(n3006), .Y(n771) );
  MXI2XL U1874 ( .A(n1658), .B(n2144), .S0(n3006), .Y(n770) );
  MXI2XL U1875 ( .A(n1659), .B(n2142), .S0(n3006), .Y(n769) );
  MXI2XL U1876 ( .A(n1660), .B(n2202), .S0(n3006), .Y(n768) );
  MXI2XL U1877 ( .A(n1661), .B(n2200), .S0(n3006), .Y(n767) );
  MXI2XL U1878 ( .A(n1662), .B(n2198), .S0(n3006), .Y(n766) );
  MXI2XL U1879 ( .A(n1663), .B(n2196), .S0(n3006), .Y(n765) );
  MXI2XL U1880 ( .A(n1664), .B(n2194), .S0(n3006), .Y(n764) );
  MXI2XL U1881 ( .A(n1665), .B(n2192), .S0(n3006), .Y(n763) );
  MXI2XL U1882 ( .A(n1666), .B(n2190), .S0(n3006), .Y(n762) );
  MXI2XL U1883 ( .A(n1667), .B(n2188), .S0(n3006), .Y(n761) );
  MXI2XL U1884 ( .A(n1668), .B(n2186), .S0(n3006), .Y(n760) );
  MXI2XL U1885 ( .A(n1669), .B(n2184), .S0(n3006), .Y(n759) );
  MXI2XL U1886 ( .A(n1670), .B(n2180), .S0(n3006), .Y(n758) );
  MXI2XL U1887 ( .A(n1671), .B(n2178), .S0(n3006), .Y(n757) );
  MXI2XL U1888 ( .A(n1672), .B(n2176), .S0(n3006), .Y(n756) );
  MXI2XL U1889 ( .A(n1673), .B(n2174), .S0(n3006), .Y(n755) );
  MXI2XL U1890 ( .A(n1674), .B(n2172), .S0(n3006), .Y(n754) );
  MXI2XL U1891 ( .A(n1675), .B(n2170), .S0(n3006), .Y(n753) );
  MXI2XL U1892 ( .A(n1676), .B(n2168), .S0(n3006), .Y(n752) );
  MXI2XL U1893 ( .A(n1677), .B(n2166), .S0(n3006), .Y(n751) );
  MXI2XL U1894 ( .A(n1678), .B(n2164), .S0(n3006), .Y(n750) );
  MXI2XL U1895 ( .A(n1679), .B(n2162), .S0(n3006), .Y(n749) );
  MXI2XL U1896 ( .A(n1680), .B(n2158), .S0(n3006), .Y(n748) );
  MXI2XL U1897 ( .A(n1681), .B(n2156), .S0(n3006), .Y(n747) );
  MXI2XL U1898 ( .A(n1682), .B(n2204), .S0(n3008), .Y(n746) );
  MXI2XL U1899 ( .A(n1683), .B(n2182), .S0(n3008), .Y(n745) );
  MXI2XL U1900 ( .A(n1684), .B(n2160), .S0(n3008), .Y(n744) );
  MXI2XL U1901 ( .A(n1685), .B(n2154), .S0(n3008), .Y(n743) );
  MXI2XL U1902 ( .A(n1686), .B(n2152), .S0(n3008), .Y(n742) );
  MXI2XL U1903 ( .A(n1687), .B(n2150), .S0(n3008), .Y(n741) );
  MXI2XL U1904 ( .A(n1688), .B(n2148), .S0(n3008), .Y(n740) );
  MXI2XL U1905 ( .A(n1689), .B(n2146), .S0(n3008), .Y(n739) );
  MXI2XL U1906 ( .A(n1690), .B(n2144), .S0(n3008), .Y(n738) );
  MXI2XL U1907 ( .A(n1691), .B(n2142), .S0(n3008), .Y(n737) );
  MXI2XL U1908 ( .A(n1692), .B(n2202), .S0(n3008), .Y(n736) );
  MXI2XL U1909 ( .A(n1693), .B(n2200), .S0(n3008), .Y(n735) );
  MXI2XL U1910 ( .A(n1694), .B(n2198), .S0(n3008), .Y(n734) );
  MXI2XL U1911 ( .A(n1695), .B(n2196), .S0(n3008), .Y(n733) );
  MXI2XL U1912 ( .A(n1696), .B(n2194), .S0(n3008), .Y(n732) );
  MXI2XL U1913 ( .A(n1697), .B(n2192), .S0(n3008), .Y(n731) );
  MXI2XL U1914 ( .A(n1698), .B(n2190), .S0(n3008), .Y(n730) );
  MXI2XL U1915 ( .A(n1699), .B(n2188), .S0(n3008), .Y(n729) );
  MXI2XL U1916 ( .A(n1700), .B(n2186), .S0(n3008), .Y(n728) );
  MXI2XL U1917 ( .A(n1701), .B(n2184), .S0(n3008), .Y(n727) );
  MXI2XL U1918 ( .A(n1702), .B(n2180), .S0(n3008), .Y(n726) );
  MXI2XL U1919 ( .A(n1703), .B(n2178), .S0(n3008), .Y(n725) );
  MXI2XL U1920 ( .A(n1704), .B(n2176), .S0(n3008), .Y(n724) );
  MXI2XL U1921 ( .A(n1705), .B(n2174), .S0(n3008), .Y(n723) );
  MXI2XL U1922 ( .A(n1706), .B(n2172), .S0(n3008), .Y(n722) );
  MXI2XL U1923 ( .A(n1707), .B(n2170), .S0(n3008), .Y(n721) );
  MXI2XL U1924 ( .A(n1708), .B(n2168), .S0(n3008), .Y(n720) );
  MXI2XL U1925 ( .A(n1709), .B(n2166), .S0(n3008), .Y(n719) );
  MXI2XL U1926 ( .A(n1710), .B(n2164), .S0(n3008), .Y(n718) );
  MXI2XL U1927 ( .A(n1711), .B(n2162), .S0(n3008), .Y(n717) );
  MXI2XL U1928 ( .A(n1712), .B(n2158), .S0(n3008), .Y(n716) );
  MXI2XL U1929 ( .A(n1713), .B(n2156), .S0(n3008), .Y(n715) );
  MXI2XL U1930 ( .A(n1714), .B(n2204), .S0(n3010), .Y(n714) );
  MXI2XL U1931 ( .A(n1715), .B(n2182), .S0(n3010), .Y(n713) );
  MXI2XL U1932 ( .A(n1716), .B(n2160), .S0(n3010), .Y(n712) );
  MXI2XL U1933 ( .A(n1717), .B(n2154), .S0(n3010), .Y(n711) );
  MXI2XL U1934 ( .A(n1718), .B(n2152), .S0(n3010), .Y(n710) );
  MXI2XL U1935 ( .A(n1719), .B(n2150), .S0(n3010), .Y(n709) );
  MXI2XL U1936 ( .A(n1720), .B(n2148), .S0(n3010), .Y(n708) );
  MXI2XL U1937 ( .A(n1721), .B(n2146), .S0(n3010), .Y(n707) );
  MXI2XL U1938 ( .A(n1722), .B(n2144), .S0(n3010), .Y(n706) );
  MXI2XL U1939 ( .A(n1723), .B(n2142), .S0(n3010), .Y(n705) );
  MXI2XL U1940 ( .A(n1724), .B(n2202), .S0(n3010), .Y(n704) );
  MXI2XL U1941 ( .A(n1725), .B(n2200), .S0(n3010), .Y(n703) );
  MXI2XL U1942 ( .A(n1726), .B(n2198), .S0(n3010), .Y(n702) );
  MXI2XL U1943 ( .A(n1727), .B(n2196), .S0(n3010), .Y(n701) );
  MXI2XL U1944 ( .A(n1728), .B(n2194), .S0(n3010), .Y(n700) );
  MXI2XL U1945 ( .A(n1729), .B(n2192), .S0(n3010), .Y(n699) );
  MXI2XL U1946 ( .A(n1730), .B(n2190), .S0(n3010), .Y(n698) );
  MXI2XL U1947 ( .A(n1731), .B(n2188), .S0(n3010), .Y(n697) );
  MXI2XL U1948 ( .A(n1732), .B(n2186), .S0(n3010), .Y(n696) );
  MXI2XL U1949 ( .A(n1733), .B(n2184), .S0(n3010), .Y(n695) );
  MXI2XL U1950 ( .A(n1734), .B(n2180), .S0(n3010), .Y(n694) );
  MXI2XL U1951 ( .A(n1735), .B(n2178), .S0(n3010), .Y(n693) );
  MXI2XL U1952 ( .A(n1736), .B(n2176), .S0(n3010), .Y(n692) );
  MXI2XL U1953 ( .A(n1737), .B(n2174), .S0(n3010), .Y(n691) );
  MXI2XL U1954 ( .A(n1738), .B(n2172), .S0(n3010), .Y(n690) );
  MXI2XL U1955 ( .A(n1739), .B(n2170), .S0(n3010), .Y(n689) );
  MXI2XL U1956 ( .A(n1740), .B(n2168), .S0(n3010), .Y(n688) );
  MXI2XL U1957 ( .A(n1741), .B(n2166), .S0(n3010), .Y(n687) );
  MXI2XL U1958 ( .A(n1742), .B(n2164), .S0(n3010), .Y(n686) );
  MXI2XL U1959 ( .A(n1743), .B(n2162), .S0(n3010), .Y(n685) );
  MXI2XL U1960 ( .A(n1744), .B(n2158), .S0(n3010), .Y(n684) );
  MXI2XL U1961 ( .A(n1745), .B(n2156), .S0(n3010), .Y(n683) );
  MXI2XL U1962 ( .A(n1746), .B(n2204), .S0(n3011), .Y(n682) );
  MXI2XL U1963 ( .A(n1747), .B(n2182), .S0(n3011), .Y(n681) );
  MXI2XL U1964 ( .A(n1748), .B(n2160), .S0(n3011), .Y(n680) );
  MXI2XL U1965 ( .A(n1749), .B(n2154), .S0(n3011), .Y(n679) );
  MXI2XL U1966 ( .A(n1750), .B(n2152), .S0(n3011), .Y(n678) );
  MXI2XL U1967 ( .A(n1751), .B(n2150), .S0(n3011), .Y(n677) );
  MXI2XL U1968 ( .A(n1752), .B(n2148), .S0(n3011), .Y(n676) );
  MXI2XL U1969 ( .A(n1753), .B(n2146), .S0(n3011), .Y(n675) );
  MXI2XL U1970 ( .A(n1754), .B(n2144), .S0(n3011), .Y(n674) );
  MXI2XL U1971 ( .A(n1755), .B(n2142), .S0(n3011), .Y(n673) );
  MXI2XL U1972 ( .A(n1756), .B(n2202), .S0(n3011), .Y(n672) );
  MXI2XL U1973 ( .A(n1757), .B(n2200), .S0(n3011), .Y(n671) );
  MXI2XL U1974 ( .A(n1758), .B(n2198), .S0(n3011), .Y(n670) );
  MXI2XL U1975 ( .A(n1759), .B(n2196), .S0(n3011), .Y(n669) );
  MXI2XL U1976 ( .A(n1760), .B(n2194), .S0(n3011), .Y(n668) );
  MXI2XL U1977 ( .A(n1761), .B(n2192), .S0(n3011), .Y(n667) );
  MXI2XL U1978 ( .A(n1762), .B(n2190), .S0(n3011), .Y(n666) );
  MXI2XL U1979 ( .A(n1763), .B(n2188), .S0(n3011), .Y(n665) );
  MXI2XL U1980 ( .A(n1764), .B(n2186), .S0(n3011), .Y(n664) );
  MXI2XL U1981 ( .A(n1765), .B(n2184), .S0(n3011), .Y(n663) );
  MXI2XL U1982 ( .A(n1766), .B(n2180), .S0(n3011), .Y(n662) );
  MXI2XL U1983 ( .A(n1767), .B(n2178), .S0(n3011), .Y(n661) );
  MXI2XL U1984 ( .A(n1768), .B(n2176), .S0(n3011), .Y(n660) );
  MXI2XL U1985 ( .A(n1769), .B(n2174), .S0(n3011), .Y(n659) );
  MXI2XL U1986 ( .A(n1770), .B(n2172), .S0(n3011), .Y(n658) );
  MXI2XL U1987 ( .A(n1771), .B(n2170), .S0(n3011), .Y(n657) );
  MXI2XL U1988 ( .A(n1772), .B(n2168), .S0(n3011), .Y(n656) );
  MXI2XL U1989 ( .A(n1773), .B(n2166), .S0(n3011), .Y(n655) );
  MXI2XL U1990 ( .A(n1774), .B(n2164), .S0(n3011), .Y(n654) );
  MXI2XL U1991 ( .A(n1775), .B(n2162), .S0(n3011), .Y(n653) );
  MXI2XL U1992 ( .A(n1776), .B(n2158), .S0(n3011), .Y(n652) );
  MXI2XL U1993 ( .A(n1777), .B(n2156), .S0(n3011), .Y(n651) );
  MXI2XL U1994 ( .A(n1778), .B(n2204), .S0(n3012), .Y(n650) );
  MXI2XL U1995 ( .A(n1779), .B(n2182), .S0(n3012), .Y(n649) );
  MXI2XL U1996 ( .A(n1780), .B(n2160), .S0(n3012), .Y(n648) );
  MXI2XL U1997 ( .A(n1781), .B(n2154), .S0(n3012), .Y(n647) );
  MXI2XL U1998 ( .A(n1782), .B(n2152), .S0(n3012), .Y(n646) );
  MXI2XL U1999 ( .A(n1783), .B(n2150), .S0(n3012), .Y(n645) );
  MXI2XL U2000 ( .A(n1784), .B(n2148), .S0(n3012), .Y(n644) );
  MXI2XL U2001 ( .A(n1785), .B(n2146), .S0(n3012), .Y(n643) );
  MXI2XL U2002 ( .A(n1786), .B(n2144), .S0(n3012), .Y(n642) );
  MXI2XL U2003 ( .A(n1787), .B(n2142), .S0(n3012), .Y(n641) );
  MXI2XL U2004 ( .A(n1788), .B(n2202), .S0(n3012), .Y(n640) );
  MXI2XL U2005 ( .A(n1789), .B(n2200), .S0(n3012), .Y(n639) );
  MXI2XL U2006 ( .A(n1790), .B(n2198), .S0(n3012), .Y(n638) );
  MXI2XL U2007 ( .A(n1791), .B(n2196), .S0(n3012), .Y(n637) );
  MXI2XL U2008 ( .A(n1792), .B(n2194), .S0(n3012), .Y(n636) );
  MXI2XL U2009 ( .A(n1793), .B(n2192), .S0(n3012), .Y(n635) );
  MXI2XL U2010 ( .A(n1794), .B(n2190), .S0(n3012), .Y(n634) );
  MXI2XL U2011 ( .A(n1795), .B(n2188), .S0(n3012), .Y(n633) );
  MXI2XL U2012 ( .A(n1796), .B(n2186), .S0(n3012), .Y(n632) );
  MXI2XL U2013 ( .A(n1797), .B(n2184), .S0(n3012), .Y(n631) );
  MXI2XL U2014 ( .A(n1798), .B(n2180), .S0(n3012), .Y(n630) );
  MXI2XL U2015 ( .A(n1799), .B(n2178), .S0(n3012), .Y(n629) );
  MXI2XL U2016 ( .A(n1800), .B(n2176), .S0(n3012), .Y(n628) );
  MXI2XL U2017 ( .A(n1801), .B(n2174), .S0(n3012), .Y(n627) );
  MXI2XL U2018 ( .A(n1802), .B(n2172), .S0(n3012), .Y(n626) );
  MXI2XL U2019 ( .A(n1803), .B(n2170), .S0(n3012), .Y(n625) );
  MXI2XL U2020 ( .A(n1804), .B(n2168), .S0(n3012), .Y(n624) );
  MXI2XL U2021 ( .A(n1805), .B(n2166), .S0(n3012), .Y(n623) );
  MXI2XL U2022 ( .A(n1806), .B(n2164), .S0(n3012), .Y(n622) );
  MXI2XL U2023 ( .A(n1807), .B(n2162), .S0(n3012), .Y(n621) );
  MXI2XL U2024 ( .A(n1808), .B(n2158), .S0(n3012), .Y(n620) );
  MXI2XL U2025 ( .A(n1809), .B(n2156), .S0(n3012), .Y(n619) );
  MXI2XL U2026 ( .A(n1810), .B(n2204), .S0(n3013), .Y(n618) );
  MXI2XL U2027 ( .A(n1811), .B(n2182), .S0(n3013), .Y(n617) );
  MXI2XL U2028 ( .A(n1812), .B(n2160), .S0(n3013), .Y(n616) );
  MXI2XL U2029 ( .A(n1813), .B(n2154), .S0(n3013), .Y(n615) );
  MXI2XL U2030 ( .A(n1814), .B(n2152), .S0(n3013), .Y(n614) );
  MXI2XL U2031 ( .A(n1815), .B(n2150), .S0(n3013), .Y(n613) );
  MXI2XL U2032 ( .A(n1816), .B(n2148), .S0(n3013), .Y(n612) );
  MXI2XL U2033 ( .A(n1817), .B(n2146), .S0(n3013), .Y(n611) );
  MXI2XL U2034 ( .A(n1818), .B(n2144), .S0(n3013), .Y(n610) );
  MXI2XL U2035 ( .A(n1819), .B(n2142), .S0(n3013), .Y(n609) );
  MXI2XL U2036 ( .A(n1820), .B(n2202), .S0(n3013), .Y(n608) );
  MXI2XL U2037 ( .A(n1821), .B(n2200), .S0(n3013), .Y(n607) );
  MXI2XL U2038 ( .A(n1822), .B(n2198), .S0(n3013), .Y(n606) );
  MXI2XL U2039 ( .A(n1823), .B(n2196), .S0(n3013), .Y(n605) );
  MXI2XL U2040 ( .A(n1824), .B(n2194), .S0(n3013), .Y(n604) );
  MXI2XL U2041 ( .A(n1825), .B(n2192), .S0(n3013), .Y(n603) );
  MXI2XL U2042 ( .A(n1826), .B(n2190), .S0(n3013), .Y(n602) );
  MXI2XL U2043 ( .A(n1827), .B(n2188), .S0(n3013), .Y(n601) );
  MXI2XL U2044 ( .A(n1828), .B(n2186), .S0(n3013), .Y(n600) );
  MXI2XL U2045 ( .A(n1829), .B(n2184), .S0(n3013), .Y(n599) );
  MXI2XL U2046 ( .A(n1830), .B(n2180), .S0(n3013), .Y(n598) );
  MXI2XL U2047 ( .A(n1831), .B(n2178), .S0(n3013), .Y(n597) );
  MXI2XL U2048 ( .A(n1832), .B(n2176), .S0(n3013), .Y(n596) );
  MXI2XL U2049 ( .A(n1833), .B(n2174), .S0(n3013), .Y(n595) );
  MXI2XL U2050 ( .A(n1834), .B(n2172), .S0(n3013), .Y(n594) );
  MXI2XL U2051 ( .A(n1835), .B(n2170), .S0(n3013), .Y(n593) );
  MXI2XL U2052 ( .A(n1836), .B(n2168), .S0(n3013), .Y(n592) );
  MXI2XL U2053 ( .A(n1837), .B(n2166), .S0(n3013), .Y(n591) );
  MXI2XL U2054 ( .A(n1838), .B(n2164), .S0(n3013), .Y(n590) );
  MXI2XL U2055 ( .A(n1839), .B(n2162), .S0(n3013), .Y(n589) );
  MXI2XL U2056 ( .A(n1840), .B(n2158), .S0(n3013), .Y(n588) );
  MXI2XL U2057 ( .A(n1841), .B(n2156), .S0(n3013), .Y(n587) );
  MXI2XL U2058 ( .A(n1842), .B(n2204), .S0(n3014), .Y(n586) );
  MXI2XL U2059 ( .A(n1843), .B(n2182), .S0(n3014), .Y(n585) );
  MXI2XL U2060 ( .A(n1844), .B(n2160), .S0(n3014), .Y(n584) );
  MXI2XL U2061 ( .A(n1845), .B(n2154), .S0(n3014), .Y(n583) );
  MXI2XL U2062 ( .A(n1846), .B(n2152), .S0(n3014), .Y(n582) );
  MXI2XL U2063 ( .A(n1847), .B(n2150), .S0(n3014), .Y(n581) );
  MXI2XL U2064 ( .A(n1848), .B(n2148), .S0(n3014), .Y(n580) );
  MXI2XL U2065 ( .A(n1849), .B(n2146), .S0(n3014), .Y(n579) );
  MXI2XL U2066 ( .A(n1850), .B(n2144), .S0(n3014), .Y(n578) );
  MXI2XL U2067 ( .A(n1851), .B(n2142), .S0(n3014), .Y(n577) );
  MXI2XL U2068 ( .A(n1852), .B(n2202), .S0(n3014), .Y(n576) );
  MXI2XL U2069 ( .A(n1853), .B(n2200), .S0(n3014), .Y(n575) );
  MXI2XL U2070 ( .A(n1854), .B(n2198), .S0(n3014), .Y(n574) );
  MXI2XL U2071 ( .A(n1855), .B(n2196), .S0(n3014), .Y(n573) );
  MXI2XL U2072 ( .A(n1856), .B(n2194), .S0(n3014), .Y(n572) );
  MXI2XL U2073 ( .A(n1857), .B(n2192), .S0(n3014), .Y(n571) );
  MXI2XL U2074 ( .A(n1858), .B(n2190), .S0(n3014), .Y(n570) );
  MXI2XL U2075 ( .A(n1859), .B(n2188), .S0(n3014), .Y(n569) );
  MXI2XL U2076 ( .A(n1860), .B(n2186), .S0(n3014), .Y(n568) );
  MXI2XL U2077 ( .A(n1861), .B(n2184), .S0(n3014), .Y(n567) );
  MXI2XL U2078 ( .A(n1862), .B(n2180), .S0(n3014), .Y(n566) );
  MXI2XL U2079 ( .A(n1863), .B(n2178), .S0(n3014), .Y(n565) );
  MXI2XL U2080 ( .A(n1864), .B(n2176), .S0(n3014), .Y(n564) );
  MXI2XL U2081 ( .A(n1865), .B(n2174), .S0(n3014), .Y(n563) );
  MXI2XL U2082 ( .A(n1866), .B(n2172), .S0(n3014), .Y(n562) );
  MXI2XL U2083 ( .A(n1867), .B(n2170), .S0(n3014), .Y(n561) );
  MXI2XL U2084 ( .A(n1868), .B(n2168), .S0(n3014), .Y(n560) );
  MXI2XL U2085 ( .A(n1869), .B(n2166), .S0(n3014), .Y(n559) );
  MXI2XL U2086 ( .A(n1870), .B(n2164), .S0(n3014), .Y(n558) );
  MXI2XL U2087 ( .A(n1871), .B(n2162), .S0(n3014), .Y(n557) );
  MXI2XL U2088 ( .A(n1872), .B(n2158), .S0(n3014), .Y(n556) );
  MXI2XL U2089 ( .A(n1873), .B(n2156), .S0(n3014), .Y(n555) );
  MXI2XL U2090 ( .A(n1874), .B(n2204), .S0(n3016), .Y(n554) );
  MXI2XL U2091 ( .A(n1875), .B(n2182), .S0(n3016), .Y(n553) );
  MXI2XL U2092 ( .A(n1876), .B(n2160), .S0(n3016), .Y(n552) );
  MXI2XL U2093 ( .A(n1877), .B(n2154), .S0(n3016), .Y(n551) );
  MXI2XL U2094 ( .A(n1878), .B(n2152), .S0(n3016), .Y(n550) );
  MXI2XL U2095 ( .A(n1879), .B(n2150), .S0(n3016), .Y(n549) );
  MXI2XL U2096 ( .A(n1880), .B(n2148), .S0(n3016), .Y(n548) );
  MXI2XL U2097 ( .A(n1881), .B(n2146), .S0(n3016), .Y(n547) );
  MXI2XL U2098 ( .A(n1882), .B(n2144), .S0(n3016), .Y(n546) );
  MXI2XL U2099 ( .A(n1883), .B(n2142), .S0(n3016), .Y(n545) );
  MXI2XL U2100 ( .A(n1884), .B(n2202), .S0(n3016), .Y(n544) );
  MXI2XL U2101 ( .A(n1885), .B(n2200), .S0(n3016), .Y(n543) );
  MXI2XL U2102 ( .A(n1886), .B(n2198), .S0(n3016), .Y(n542) );
  MXI2XL U2103 ( .A(n1887), .B(n2196), .S0(n3016), .Y(n541) );
  MXI2XL U2104 ( .A(n1888), .B(n2194), .S0(n3016), .Y(n540) );
  MXI2XL U2105 ( .A(n1889), .B(n2192), .S0(n3016), .Y(n539) );
  MXI2XL U2106 ( .A(n1890), .B(n2190), .S0(n3016), .Y(n538) );
  MXI2XL U2107 ( .A(n1891), .B(n2188), .S0(n3016), .Y(n537) );
  MXI2XL U2108 ( .A(n1892), .B(n2186), .S0(n3016), .Y(n536) );
  MXI2XL U2109 ( .A(n1893), .B(n2184), .S0(n3016), .Y(n535) );
  MXI2XL U2110 ( .A(n1894), .B(n2180), .S0(n3016), .Y(n534) );
  MXI2XL U2111 ( .A(n1895), .B(n2178), .S0(n3016), .Y(n533) );
  MXI2XL U2112 ( .A(n1896), .B(n2176), .S0(n3016), .Y(n532) );
  MXI2XL U2113 ( .A(n1897), .B(n2174), .S0(n3016), .Y(n531) );
  MXI2XL U2114 ( .A(n1898), .B(n2172), .S0(n3016), .Y(n530) );
  MXI2XL U2115 ( .A(n1899), .B(n2170), .S0(n3016), .Y(n529) );
  MXI2XL U2116 ( .A(n1900), .B(n2168), .S0(n3016), .Y(n528) );
  MXI2XL U2117 ( .A(n1901), .B(n2166), .S0(n3016), .Y(n527) );
  MXI2XL U2118 ( .A(n1902), .B(n2164), .S0(n3016), .Y(n526) );
  MXI2XL U2119 ( .A(n1903), .B(n2162), .S0(n3016), .Y(n525) );
  MXI2XL U2120 ( .A(n1904), .B(n2158), .S0(n3016), .Y(n524) );
  MXI2XL U2121 ( .A(n1905), .B(n2156), .S0(n3016), .Y(n523) );
  MXI2XL U2122 ( .A(n1906), .B(n2204), .S0(n3018), .Y(n522) );
  MXI2XL U2123 ( .A(n1907), .B(n2182), .S0(n3018), .Y(n521) );
  MXI2XL U2124 ( .A(n1908), .B(n2160), .S0(n3018), .Y(n520) );
  MXI2XL U2125 ( .A(n1909), .B(n2154), .S0(n3018), .Y(n519) );
  MXI2XL U2126 ( .A(n1910), .B(n2152), .S0(n3018), .Y(n518) );
  MXI2XL U2127 ( .A(n1911), .B(n2150), .S0(n3018), .Y(n517) );
  MXI2XL U2128 ( .A(n1912), .B(n2148), .S0(n3018), .Y(n516) );
  MXI2XL U2129 ( .A(n1913), .B(n2146), .S0(n3018), .Y(n515) );
  MXI2XL U2130 ( .A(n1914), .B(n2144), .S0(n3018), .Y(n514) );
  MXI2XL U2131 ( .A(n1915), .B(n2142), .S0(n3018), .Y(n513) );
  MXI2XL U2132 ( .A(n1916), .B(n2202), .S0(n3018), .Y(n512) );
  MXI2XL U2133 ( .A(n1917), .B(n2200), .S0(n3018), .Y(n511) );
  MXI2XL U2134 ( .A(n1918), .B(n2198), .S0(n3018), .Y(n510) );
  MXI2XL U2135 ( .A(n1919), .B(n2196), .S0(n3018), .Y(n509) );
  MXI2XL U2136 ( .A(n1920), .B(n2194), .S0(n3018), .Y(n508) );
  MXI2XL U2137 ( .A(n1921), .B(n2192), .S0(n3018), .Y(n507) );
  MXI2XL U2138 ( .A(n1922), .B(n2190), .S0(n3018), .Y(n506) );
  MXI2XL U2139 ( .A(n1923), .B(n2188), .S0(n3018), .Y(n505) );
  MXI2XL U2140 ( .A(n1924), .B(n2186), .S0(n3018), .Y(n504) );
  MXI2XL U2141 ( .A(n1925), .B(n2184), .S0(n3018), .Y(n503) );
  MXI2XL U2142 ( .A(n1926), .B(n2180), .S0(n3018), .Y(n502) );
  MXI2XL U2143 ( .A(n1927), .B(n2178), .S0(n3018), .Y(n501) );
  MXI2XL U2144 ( .A(n1928), .B(n2176), .S0(n3018), .Y(n500) );
  MXI2XL U2145 ( .A(n1929), .B(n2174), .S0(n3018), .Y(n499) );
  MXI2XL U2146 ( .A(n1930), .B(n2172), .S0(n3018), .Y(n498) );
  MXI2XL U2147 ( .A(n1931), .B(n2170), .S0(n3018), .Y(n497) );
  MXI2XL U2148 ( .A(n1932), .B(n2168), .S0(n3018), .Y(n496) );
  MXI2XL U2149 ( .A(n1933), .B(n2166), .S0(n3018), .Y(n495) );
  MXI2XL U2150 ( .A(n1934), .B(n2164), .S0(n3018), .Y(n494) );
  MXI2XL U2151 ( .A(n1935), .B(n2162), .S0(n3018), .Y(n493) );
  MXI2XL U2152 ( .A(n1936), .B(n2158), .S0(n3018), .Y(n492) );
  MXI2XL U2153 ( .A(n1937), .B(n2156), .S0(n3018), .Y(n491) );
  MXI2XL U2154 ( .A(n1938), .B(n2204), .S0(n3019), .Y(n490) );
  MXI2XL U2155 ( .A(n1939), .B(n2182), .S0(n3019), .Y(n489) );
  MXI2XL U2156 ( .A(n1940), .B(n2160), .S0(n3019), .Y(n488) );
  MXI2XL U2157 ( .A(n1941), .B(n2154), .S0(n3019), .Y(n487) );
  MXI2XL U2158 ( .A(n1942), .B(n2152), .S0(n3019), .Y(n486) );
  MXI2XL U2159 ( .A(n1943), .B(n2150), .S0(n3019), .Y(n485) );
  MXI2XL U2160 ( .A(n1944), .B(n2148), .S0(n3019), .Y(n484) );
  MXI2XL U2161 ( .A(n1945), .B(n2146), .S0(n3019), .Y(n483) );
  MXI2XL U2162 ( .A(n1946), .B(n2144), .S0(n3019), .Y(n482) );
  MXI2XL U2163 ( .A(n1947), .B(n2142), .S0(n3019), .Y(n481) );
  MXI2XL U2164 ( .A(n1948), .B(n2202), .S0(n3019), .Y(n480) );
  MXI2XL U2165 ( .A(n1949), .B(n2200), .S0(n3019), .Y(n479) );
  MXI2XL U2166 ( .A(n1950), .B(n2198), .S0(n3019), .Y(n478) );
  MXI2XL U2167 ( .A(n1951), .B(n2196), .S0(n3019), .Y(n477) );
  MXI2XL U2168 ( .A(n1952), .B(n2194), .S0(n3019), .Y(n476) );
  MXI2XL U2169 ( .A(n1953), .B(n2192), .S0(n3019), .Y(n475) );
  MXI2XL U2170 ( .A(n1954), .B(n2190), .S0(n3019), .Y(n474) );
  MXI2XL U2171 ( .A(n1955), .B(n2188), .S0(n3019), .Y(n473) );
  MXI2XL U2172 ( .A(n1956), .B(n2186), .S0(n3019), .Y(n472) );
  MXI2XL U2173 ( .A(n1957), .B(n2184), .S0(n3019), .Y(n471) );
  MXI2XL U2174 ( .A(n1958), .B(n2180), .S0(n3019), .Y(n470) );
  MXI2XL U2175 ( .A(n1959), .B(n2178), .S0(n3019), .Y(n469) );
  MXI2XL U2176 ( .A(n1960), .B(n2176), .S0(n3019), .Y(n468) );
  MXI2XL U2177 ( .A(n1961), .B(n2174), .S0(n3019), .Y(n467) );
  MXI2XL U2178 ( .A(n1962), .B(n2172), .S0(n3019), .Y(n466) );
  MXI2XL U2179 ( .A(n1963), .B(n2170), .S0(n3019), .Y(n465) );
  MXI2XL U2180 ( .A(n1964), .B(n2168), .S0(n3019), .Y(n464) );
  MXI2XL U2181 ( .A(n1965), .B(n2166), .S0(n3019), .Y(n463) );
  MXI2XL U2182 ( .A(n1966), .B(n2164), .S0(n3019), .Y(n462) );
  MXI2XL U2183 ( .A(n1967), .B(n2162), .S0(n3019), .Y(n461) );
  MXI2XL U2184 ( .A(n1968), .B(n2158), .S0(n3019), .Y(n460) );
  MXI2XL U2185 ( .A(n1969), .B(n2156), .S0(n3019), .Y(n459) );
  MXI2XL U2186 ( .A(n1970), .B(n2204), .S0(n3020), .Y(n458) );
  MXI2XL U2187 ( .A(n1971), .B(n2182), .S0(n3020), .Y(n457) );
  MXI2XL U2188 ( .A(n1972), .B(n2160), .S0(n3020), .Y(n456) );
  MXI2XL U2189 ( .A(n1973), .B(n2154), .S0(n3020), .Y(n455) );
  MXI2XL U2190 ( .A(n1974), .B(n2152), .S0(n3020), .Y(n454) );
  MXI2XL U2191 ( .A(n1975), .B(n2150), .S0(n3020), .Y(n453) );
  MXI2XL U2192 ( .A(n1976), .B(n2148), .S0(n3020), .Y(n452) );
  MXI2XL U2193 ( .A(n1977), .B(n2146), .S0(n3020), .Y(n451) );
  MXI2XL U2194 ( .A(n1978), .B(n2144), .S0(n3020), .Y(n450) );
  MXI2XL U2195 ( .A(n1979), .B(n2142), .S0(n3020), .Y(n449) );
  MXI2XL U2196 ( .A(n1980), .B(n2202), .S0(n3020), .Y(n448) );
  MXI2XL U2197 ( .A(n1981), .B(n2200), .S0(n3020), .Y(n447) );
  MXI2XL U2198 ( .A(n1982), .B(n2198), .S0(n3020), .Y(n446) );
  MXI2XL U2199 ( .A(n1983), .B(n2196), .S0(n3020), .Y(n445) );
  MXI2XL U2200 ( .A(n1984), .B(n2194), .S0(n3020), .Y(n444) );
  MXI2XL U2201 ( .A(n1985), .B(n2192), .S0(n3020), .Y(n443) );
  MXI2XL U2202 ( .A(n1986), .B(n2190), .S0(n3020), .Y(n442) );
  MXI2XL U2203 ( .A(n1987), .B(n2188), .S0(n3020), .Y(n441) );
  MXI2XL U2204 ( .A(n1988), .B(n2186), .S0(n3020), .Y(n440) );
  MXI2XL U2205 ( .A(n1989), .B(n2184), .S0(n3020), .Y(n439) );
  MXI2XL U2206 ( .A(n1990), .B(n2180), .S0(n3020), .Y(n438) );
  MXI2XL U2207 ( .A(n1991), .B(n2178), .S0(n3020), .Y(n437) );
  MXI2XL U2208 ( .A(n1992), .B(n2176), .S0(n3020), .Y(n436) );
  MXI2XL U2209 ( .A(n1993), .B(n2174), .S0(n3020), .Y(n435) );
  MXI2XL U2210 ( .A(n1994), .B(n2172), .S0(n3020), .Y(n434) );
  MXI2XL U2211 ( .A(n1995), .B(n2170), .S0(n3020), .Y(n433) );
  MXI2XL U2212 ( .A(n1996), .B(n2168), .S0(n3020), .Y(n432) );
  MXI2XL U2213 ( .A(n1997), .B(n2166), .S0(n3020), .Y(n431) );
  MXI2XL U2214 ( .A(n1998), .B(n2164), .S0(n3020), .Y(n430) );
  MXI2XL U2215 ( .A(n1999), .B(n2162), .S0(n3020), .Y(n429) );
  MXI2XL U2216 ( .A(n2000), .B(n2158), .S0(n3020), .Y(n428) );
  MXI2XL U2217 ( .A(n2001), .B(n2156), .S0(n3020), .Y(n427) );
  MXI2XL U2218 ( .A(n2002), .B(n2204), .S0(n3021), .Y(n426) );
  MXI2XL U2219 ( .A(n2003), .B(n2182), .S0(n3021), .Y(n425) );
  MXI2XL U2220 ( .A(n2004), .B(n2160), .S0(n3021), .Y(n424) );
  MXI2XL U2221 ( .A(n2005), .B(n2154), .S0(n3021), .Y(n423) );
  MXI2XL U2222 ( .A(n2006), .B(n2152), .S0(n3021), .Y(n422) );
  MXI2XL U2223 ( .A(n2007), .B(n2150), .S0(n3021), .Y(n421) );
  MXI2XL U2224 ( .A(n2008), .B(n2148), .S0(n3021), .Y(n420) );
  MXI2XL U2225 ( .A(n2009), .B(n2146), .S0(n3021), .Y(n419) );
  MXI2XL U2226 ( .A(n2010), .B(n2144), .S0(n3021), .Y(n418) );
  MXI2XL U2227 ( .A(n2011), .B(n2142), .S0(n3021), .Y(n417) );
  MXI2XL U2228 ( .A(n2012), .B(n2202), .S0(n3021), .Y(n416) );
  MXI2XL U2229 ( .A(n2013), .B(n2200), .S0(n3021), .Y(n415) );
  MXI2XL U2230 ( .A(n2014), .B(n2198), .S0(n3021), .Y(n414) );
  MXI2XL U2231 ( .A(n2015), .B(n2196), .S0(n3021), .Y(n413) );
  MXI2XL U2232 ( .A(n2016), .B(n2194), .S0(n3021), .Y(n412) );
  MXI2XL U2233 ( .A(n2017), .B(n2192), .S0(n3021), .Y(n411) );
  MXI2XL U2234 ( .A(n2018), .B(n2190), .S0(n3021), .Y(n410) );
  MXI2XL U2235 ( .A(n2019), .B(n2188), .S0(n3021), .Y(n409) );
  MXI2XL U2236 ( .A(n2020), .B(n2186), .S0(n3021), .Y(n408) );
  MXI2XL U2237 ( .A(n2021), .B(n2184), .S0(n3021), .Y(n407) );
  MXI2XL U2238 ( .A(n2022), .B(n2180), .S0(n3021), .Y(n406) );
  MXI2XL U2239 ( .A(n2023), .B(n2178), .S0(n3021), .Y(n405) );
  MXI2XL U2240 ( .A(n2024), .B(n2176), .S0(n3021), .Y(n404) );
  MXI2XL U2241 ( .A(n2025), .B(n2174), .S0(n3021), .Y(n403) );
  MXI2XL U2242 ( .A(n2026), .B(n2172), .S0(n3021), .Y(n402) );
  MXI2XL U2243 ( .A(n2027), .B(n2170), .S0(n3021), .Y(n401) );
  MXI2XL U2244 ( .A(n2028), .B(n2168), .S0(n3021), .Y(n400) );
  MXI2XL U2245 ( .A(n2029), .B(n2166), .S0(n3021), .Y(n399) );
  MXI2XL U2246 ( .A(n2030), .B(n2164), .S0(n3021), .Y(n398) );
  MXI2XL U2247 ( .A(n2031), .B(n2162), .S0(n3021), .Y(n397) );
  MXI2XL U2248 ( .A(n2032), .B(n2158), .S0(n3021), .Y(n396) );
  MXI2XL U2249 ( .A(n2033), .B(n2156), .S0(n3021), .Y(n395) );
  MXI2XL U2250 ( .A(n2034), .B(n2204), .S0(n3022), .Y(n394) );
  MXI2XL U2251 ( .A(n2035), .B(n2182), .S0(n3022), .Y(n393) );
  MXI2XL U2252 ( .A(n2036), .B(n2160), .S0(n3022), .Y(n392) );
  MXI2XL U2253 ( .A(n2037), .B(n2154), .S0(n3022), .Y(n391) );
  MXI2XL U2254 ( .A(n2038), .B(n2152), .S0(n3022), .Y(n390) );
  MXI2XL U2255 ( .A(n2039), .B(n2150), .S0(n3022), .Y(n389) );
  MXI2XL U2256 ( .A(n2040), .B(n2148), .S0(n3022), .Y(n388) );
  MXI2XL U2257 ( .A(n2041), .B(n2146), .S0(n3022), .Y(n387) );
  MXI2XL U2258 ( .A(n2042), .B(n2144), .S0(n3022), .Y(n386) );
  MXI2XL U2259 ( .A(n2043), .B(n2142), .S0(n3022), .Y(n385) );
  MXI2XL U2260 ( .A(n2044), .B(n2202), .S0(n3022), .Y(n384) );
  MXI2XL U2261 ( .A(n2045), .B(n2200), .S0(n3022), .Y(n383) );
  MXI2XL U2262 ( .A(n2046), .B(n2198), .S0(n3022), .Y(n382) );
  MXI2XL U2263 ( .A(n2047), .B(n2196), .S0(n3022), .Y(n381) );
  MXI2XL U2264 ( .A(n2048), .B(n2194), .S0(n3022), .Y(n380) );
  MXI2XL U2265 ( .A(n2049), .B(n2192), .S0(n3022), .Y(n379) );
  MXI2XL U2266 ( .A(n2050), .B(n2190), .S0(n3022), .Y(n378) );
  MXI2XL U2267 ( .A(n2051), .B(n2188), .S0(n3022), .Y(n377) );
  MXI2XL U2268 ( .A(n2052), .B(n2186), .S0(n3022), .Y(n376) );
  MXI2XL U2269 ( .A(n2053), .B(n2184), .S0(n3022), .Y(n375) );
  MXI2XL U2270 ( .A(n2054), .B(n2180), .S0(n3022), .Y(n374) );
  MXI2XL U2271 ( .A(n2055), .B(n2178), .S0(n3022), .Y(n373) );
  MXI2XL U2272 ( .A(n2056), .B(n2176), .S0(n3022), .Y(n372) );
  MXI2XL U2273 ( .A(n2057), .B(n2174), .S0(n3022), .Y(n371) );
  MXI2XL U2274 ( .A(n2058), .B(n2172), .S0(n3022), .Y(n370) );
  MXI2XL U2275 ( .A(n2059), .B(n2170), .S0(n3022), .Y(n369) );
  MXI2XL U2276 ( .A(n2060), .B(n2168), .S0(n3022), .Y(n368) );
  MXI2XL U2277 ( .A(n2061), .B(n2166), .S0(n3022), .Y(n367) );
  MXI2XL U2278 ( .A(n2062), .B(n2164), .S0(n3022), .Y(n366) );
  MXI2XL U2279 ( .A(n2063), .B(n2162), .S0(n3022), .Y(n365) );
  MXI2XL U2280 ( .A(n2064), .B(n2158), .S0(n3022), .Y(n364) );
  MXI2XL U2281 ( .A(n2065), .B(n2156), .S0(n3022), .Y(n363) );
  MXI2XL U2282 ( .A(n2066), .B(n2204), .S0(n3023), .Y(n362) );
  MXI2XL U2283 ( .A(n2067), .B(n2182), .S0(n3023), .Y(n361) );
  MXI2XL U2284 ( .A(n2068), .B(n2160), .S0(n3023), .Y(n360) );
  MXI2XL U2285 ( .A(n2069), .B(n2154), .S0(n3023), .Y(n359) );
  MXI2XL U2286 ( .A(n2070), .B(n2152), .S0(n3023), .Y(n358) );
  MXI2XL U2287 ( .A(n2071), .B(n2150), .S0(n3023), .Y(n357) );
  MXI2XL U2288 ( .A(n2072), .B(n2148), .S0(n3023), .Y(n356) );
  MXI2XL U2289 ( .A(n2073), .B(n2146), .S0(n3023), .Y(n355) );
  MXI2XL U2290 ( .A(n2074), .B(n2144), .S0(n3023), .Y(n354) );
  MXI2XL U2291 ( .A(n2075), .B(n2142), .S0(n3023), .Y(n353) );
  MXI2XL U2292 ( .A(n2076), .B(n2202), .S0(n3023), .Y(n352) );
  MXI2XL U2293 ( .A(n2077), .B(n2200), .S0(n3023), .Y(n351) );
  MXI2XL U2294 ( .A(n2078), .B(n2198), .S0(n3023), .Y(n350) );
  MXI2XL U2295 ( .A(n2079), .B(n2196), .S0(n3023), .Y(n349) );
  MXI2XL U2296 ( .A(n2080), .B(n2194), .S0(n3023), .Y(n348) );
  MXI2XL U2297 ( .A(n2081), .B(n2192), .S0(n3023), .Y(n347) );
  MXI2XL U2298 ( .A(n2082), .B(n2190), .S0(n3023), .Y(n346) );
  MXI2XL U2299 ( .A(n2083), .B(n2188), .S0(n3023), .Y(n345) );
  MXI2XL U2300 ( .A(n2084), .B(n2186), .S0(n3023), .Y(n344) );
  MXI2XL U2301 ( .A(n2085), .B(n2184), .S0(n3023), .Y(n343) );
  MXI2XL U2302 ( .A(n2086), .B(n2180), .S0(n3023), .Y(n342) );
  MXI2XL U2303 ( .A(n2087), .B(n2178), .S0(n3023), .Y(n341) );
  MXI2XL U2304 ( .A(n2088), .B(n2176), .S0(n3023), .Y(n340) );
  MXI2XL U2305 ( .A(n2089), .B(n2174), .S0(n3023), .Y(n339) );
  MXI2XL U2306 ( .A(n2090), .B(n2172), .S0(n3023), .Y(n338) );
  MXI2XL U2307 ( .A(n2091), .B(n2170), .S0(n3023), .Y(n337) );
  MXI2XL U2308 ( .A(n2092), .B(n2168), .S0(n3023), .Y(n336) );
  MXI2XL U2309 ( .A(n2093), .B(n2166), .S0(n3023), .Y(n335) );
  MXI2XL U2310 ( .A(n2094), .B(n2164), .S0(n3023), .Y(n334) );
  MXI2XL U2311 ( .A(n2095), .B(n2162), .S0(n3023), .Y(n333) );
  MXI2XL U2312 ( .A(n2096), .B(n2158), .S0(n3023), .Y(n332) );
  MXI2XL U2313 ( .A(n2097), .B(n2156), .S0(n3023), .Y(n331) );
  MXI2XL U2314 ( .A(n2098), .B(n2204), .S0(n3024), .Y(n330) );
  MXI2XL U2315 ( .A(n2099), .B(n2182), .S0(n3024), .Y(n329) );
  MXI2XL U2316 ( .A(n2100), .B(n2160), .S0(n3024), .Y(n328) );
  MXI2XL U2317 ( .A(n2101), .B(n2154), .S0(n3024), .Y(n327) );
  MXI2XL U2318 ( .A(n2102), .B(n2152), .S0(n3024), .Y(n326) );
  MXI2XL U2319 ( .A(n2103), .B(n2150), .S0(n3024), .Y(n325) );
  MXI2XL U2320 ( .A(n2104), .B(n2148), .S0(n3024), .Y(n324) );
  MXI2XL U2321 ( .A(n2105), .B(n2146), .S0(n3024), .Y(n323) );
  MXI2XL U2322 ( .A(n2106), .B(n2144), .S0(n3024), .Y(n322) );
  MXI2XL U2323 ( .A(n2107), .B(n2142), .S0(n3024), .Y(n321) );
  MXI2XL U2324 ( .A(n2108), .B(n2202), .S0(n3024), .Y(n320) );
  MXI2XL U2325 ( .A(n2109), .B(n2200), .S0(n3024), .Y(n319) );
  MXI2XL U2326 ( .A(n2110), .B(n2198), .S0(n3024), .Y(n318) );
  MXI2XL U2327 ( .A(n2111), .B(n2196), .S0(n3024), .Y(n317) );
  MXI2XL U2328 ( .A(n2112), .B(n2194), .S0(n3024), .Y(n316) );
  MXI2XL U2329 ( .A(n2113), .B(n2192), .S0(n3024), .Y(n315) );
  MXI2XL U2330 ( .A(n2114), .B(n2190), .S0(n3024), .Y(n314) );
  MXI2XL U2331 ( .A(n2115), .B(n2188), .S0(n3024), .Y(n313) );
  MXI2XL U2332 ( .A(n2116), .B(n2186), .S0(n3024), .Y(n312) );
  MXI2XL U2333 ( .A(n2117), .B(n2184), .S0(n3024), .Y(n311) );
  MXI2XL U2334 ( .A(n2118), .B(n2180), .S0(n3024), .Y(n310) );
  MXI2XL U2335 ( .A(n2119), .B(n2178), .S0(n3024), .Y(n309) );
  MXI2XL U2336 ( .A(n2120), .B(n2176), .S0(n3024), .Y(n308) );
  MXI2XL U2337 ( .A(n2121), .B(n2174), .S0(n3024), .Y(n307) );
  MXI2XL U2338 ( .A(n2122), .B(n2172), .S0(n3024), .Y(n306) );
  MXI2XL U2339 ( .A(n2123), .B(n2170), .S0(n3024), .Y(n305) );
  MXI2XL U2340 ( .A(n2124), .B(n2168), .S0(n3024), .Y(n304) );
  MXI2XL U2341 ( .A(n2125), .B(n2166), .S0(n3024), .Y(n303) );
  MXI2XL U2342 ( .A(n2126), .B(n2164), .S0(n3024), .Y(n302) );
  MXI2XL U2343 ( .A(n2127), .B(n2162), .S0(n3024), .Y(n301) );
  MXI2XL U2344 ( .A(n2128), .B(n2158), .S0(n3024), .Y(n300) );
  MXI2XL U2345 ( .A(n2129), .B(n2156), .S0(n3024), .Y(n299) );
  MX2XL U2346 ( .A(read_data1[19]), .B(aluresult[19]), .S0(Foward_C), .Y(
        after_C_MUX[19]) );
  MX2XL U2347 ( .A(read_data2[19]), .B(aluresult[19]), .S0(Foward_D), .Y(
        after_D_MUX[19]) );
  MX2XL U2348 ( .A(read_data1[23]), .B(aluresult[23]), .S0(Foward_C), .Y(
        after_C_MUX[23]) );
  MX2XL U2349 ( .A(read_data2[23]), .B(aluresult[23]), .S0(Foward_D), .Y(
        after_D_MUX[23]) );
  MX2XL U2350 ( .A(read_data1[15]), .B(aluresult[15]), .S0(Foward_C), .Y(
        after_C_MUX[15]) );
  MX2XL U2351 ( .A(read_data2[15]), .B(aluresult[15]), .S0(Foward_D), .Y(
        after_D_MUX[15]) );
  MX2XL U2352 ( .A(read_data1[27]), .B(aluresult[27]), .S0(Foward_C), .Y(
        after_C_MUX[27]) );
  MX2XL U2353 ( .A(read_data2[27]), .B(aluresult[27]), .S0(Foward_D), .Y(
        after_D_MUX[27]) );
  MX2XL U2354 ( .A(read_data1[3]), .B(aluresult[3]), .S0(Foward_C), .Y(
        after_C_MUX[3]) );
  MX2XL U2355 ( .A(read_data2[3]), .B(aluresult[3]), .S0(Foward_D), .Y(
        after_D_MUX[3]) );
  MX2XL U2356 ( .A(read_data1[21]), .B(aluresult[21]), .S0(Foward_C), .Y(
        after_C_MUX[21]) );
  MX2XL U2357 ( .A(read_data2[21]), .B(aluresult[21]), .S0(Foward_D), .Y(
        after_D_MUX[21]) );
  MX2XL U2358 ( .A(read_data1[25]), .B(aluresult[25]), .S0(Foward_C), .Y(
        after_C_MUX[25]) );
  MX2XL U2359 ( .A(read_data2[25]), .B(aluresult[25]), .S0(Foward_D), .Y(
        after_D_MUX[25]) );
  MX2XL U2360 ( .A(read_data1[17]), .B(aluresult[17]), .S0(Foward_C), .Y(
        after_C_MUX[17]) );
  MX2XL U2361 ( .A(read_data2[17]), .B(aluresult[17]), .S0(Foward_D), .Y(
        after_D_MUX[17]) );
  MX2XL U2362 ( .A(read_data1[20]), .B(aluresult[20]), .S0(Foward_C), .Y(
        after_C_MUX[20]) );
  MX2XL U2363 ( .A(read_data2[20]), .B(aluresult[20]), .S0(Foward_D), .Y(
        after_D_MUX[20]) );
  MX2XL U2364 ( .A(read_data1[24]), .B(aluresult[24]), .S0(Foward_C), .Y(
        after_C_MUX[24]) );
  MX2XL U2365 ( .A(read_data2[24]), .B(aluresult[24]), .S0(Foward_D), .Y(
        after_D_MUX[24]) );
  MX2XL U2366 ( .A(read_data1[16]), .B(aluresult[16]), .S0(Foward_C), .Y(
        after_C_MUX[16]) );
  MX2XL U2367 ( .A(read_data2[16]), .B(aluresult[16]), .S0(Foward_D), .Y(
        after_D_MUX[16]) );
  MX2XL U2368 ( .A(read_data1[22]), .B(aluresult[22]), .S0(Foward_C), .Y(
        after_C_MUX[22]) );
  MX2XL U2369 ( .A(read_data2[22]), .B(aluresult[22]), .S0(Foward_D), .Y(
        after_D_MUX[22]) );
  MX2XL U2370 ( .A(read_data1[26]), .B(aluresult[26]), .S0(Foward_C), .Y(
        after_C_MUX[26]) );
  MX2XL U2371 ( .A(read_data2[26]), .B(aluresult[26]), .S0(Foward_D), .Y(
        after_D_MUX[26]) );
  MX2XL U2372 ( .A(read_data1[18]), .B(aluresult[18]), .S0(Foward_C), .Y(
        after_C_MUX[18]) );
  MX2XL U2373 ( .A(read_data2[18]), .B(aluresult[18]), .S0(Foward_D), .Y(
        after_D_MUX[18]) );
  NOR2BXL U2374 ( .AN(\EX[3] ), .B(n3116), .Y(EX_after_detect[3]) );
  MX2XL U2375 ( .A(read_data1[10]), .B(aluresult[10]), .S0(Foward_C), .Y(
        after_C_MUX[10]) );
  MX2XL U2376 ( .A(read_data2[10]), .B(aluresult[10]), .S0(Foward_D), .Y(
        after_D_MUX[10]) );
  MX2XL U2377 ( .A(read_data1[14]), .B(aluresult[14]), .S0(Foward_C), .Y(
        after_C_MUX[14]) );
  MX2XL U2378 ( .A(read_data2[14]), .B(aluresult[14]), .S0(Foward_D), .Y(
        after_D_MUX[14]) );
  MX2XL U2379 ( .A(read_data1[8]), .B(aluresult[8]), .S0(Foward_C), .Y(
        after_C_MUX[8]) );
  MX2XL U2380 ( .A(read_data2[8]), .B(aluresult[8]), .S0(Foward_D), .Y(
        after_D_MUX[8]) );
  MX2XL U2381 ( .A(read_data1[12]), .B(aluresult[12]), .S0(Foward_C), .Y(
        after_C_MUX[12]) );
  MX2XL U2382 ( .A(read_data2[12]), .B(aluresult[12]), .S0(Foward_D), .Y(
        after_D_MUX[12]) );
  MX2XL U2383 ( .A(read_data1[9]), .B(aluresult[9]), .S0(Foward_C), .Y(
        after_C_MUX[9]) );
  MX2XL U2384 ( .A(read_data2[9]), .B(aluresult[9]), .S0(Foward_D), .Y(
        after_D_MUX[9]) );
  MX2XL U2385 ( .A(read_data1[13]), .B(aluresult[13]), .S0(Foward_C), .Y(
        after_C_MUX[13]) );
  MX2XL U2386 ( .A(read_data2[13]), .B(aluresult[13]), .S0(Foward_D), .Y(
        after_D_MUX[13]) );
  MX2XL U2387 ( .A(read_data1[7]), .B(aluresult[7]), .S0(Foward_C), .Y(
        after_C_MUX[7]) );
  MX2XL U2388 ( .A(read_data2[7]), .B(aluresult[7]), .S0(Foward_D), .Y(
        after_D_MUX[7]) );
  MX2XL U2389 ( .A(read_data1[11]), .B(aluresult[11]), .S0(Foward_C), .Y(
        after_C_MUX[11]) );
  MX2XL U2390 ( .A(read_data2[11]), .B(aluresult[11]), .S0(Foward_D), .Y(
        after_D_MUX[11]) );
  NOR2BXL U2391 ( .AN(ALUOp[2]), .B(n3116), .Y(EX_after_detect[2]) );
  NOR2BXL U2392 ( .AN(M[1]), .B(n3116), .Y(MEM_after_detect[1]) );
  MX2XL U2393 ( .A(read_data2[29]), .B(aluresult[29]), .S0(Foward_D), .Y(
        after_D_MUX[29]) );
  MX2XL U2394 ( .A(read_data2[28]), .B(aluresult[28]), .S0(Foward_D), .Y(
        after_D_MUX[28]) );
  MX2XL U2395 ( .A(read_data2[30]), .B(aluresult[30]), .S0(Foward_D), .Y(
        after_D_MUX[30]) );
  MX2XL U2396 ( .A(read_data2[5]), .B(aluresult[5]), .S0(Foward_D), .Y(
        after_D_MUX[5]) );
  MX2XL U2397 ( .A(read_data2[4]), .B(aluresult[4]), .S0(Foward_D), .Y(
        after_D_MUX[4]) );
  MX2XL U2398 ( .A(read_data2[6]), .B(aluresult[6]), .S0(Foward_D), .Y(
        after_D_MUX[6]) );
  MX2XL U2399 ( .A(read_data2[31]), .B(aluresult[31]), .S0(Foward_D), .Y(
        after_D_MUX[31]) );
  MX2XL U2400 ( .A(read_data2[2]), .B(aluresult[2]), .S0(Foward_D), .Y(
        after_D_MUX[2]) );
  MX2XL U2401 ( .A(read_data2[1]), .B(aluresult[1]), .S0(Foward_D), .Y(
        after_D_MUX[1]) );
  MX2XL U2402 ( .A(read_data2[0]), .B(aluresult[0]), .S0(Foward_D), .Y(
        after_D_MUX[0]) );
  MX2XL U2403 ( .A(read_data1[2]), .B(aluresult[2]), .S0(Foward_C), .Y(
        after_C_MUX[2]) );
  MX2XL U2404 ( .A(read_data1[1]), .B(aluresult[1]), .S0(Foward_C), .Y(
        after_C_MUX[1]) );
  MX2XL U2405 ( .A(read_data1[0]), .B(aluresult[0]), .S0(Foward_C), .Y(
        after_C_MUX[0]) );
  MX2XL U2406 ( .A(read_data1[29]), .B(aluresult[29]), .S0(Foward_C), .Y(
        after_C_MUX[29]) );
  MX2XL U2407 ( .A(read_data1[28]), .B(aluresult[28]), .S0(Foward_C), .Y(
        after_C_MUX[28]) );
  MX2XL U2408 ( .A(read_data1[30]), .B(aluresult[30]), .S0(Foward_C), .Y(
        after_C_MUX[30]) );
  MX2XL U2409 ( .A(read_data1[5]), .B(aluresult[5]), .S0(Foward_C), .Y(
        after_C_MUX[5]) );
  MX2XL U2410 ( .A(read_data1[4]), .B(aluresult[4]), .S0(Foward_C), .Y(
        after_C_MUX[4]) );
  MX2XL U2411 ( .A(read_data1[6]), .B(aluresult[6]), .S0(Foward_C), .Y(
        after_C_MUX[6]) );
  MX2XL U2412 ( .A(read_data1[31]), .B(aluresult[31]), .S0(Foward_C), .Y(
        after_C_MUX[31]) );
  AOI2BB2XL U2413 ( .B0(EX_data1[26]), .B1(n2137), .A0N(n2168), .A1N(n2134), 
        .Y(n3146) );
  AOI2BB2XL U2414 ( .B0(EX_data1[27]), .B1(n2137), .A0N(n2166), .A1N(n2134), 
        .Y(n3144) );
  AOI2BB2XL U2415 ( .B0(EX_data1[9]), .B1(n2137), .A0N(n2142), .A1N(n2134), 
        .Y(n3119) );
  AOI2BB2XL U2416 ( .B0(EX_data1[19]), .B1(n2137), .A0N(n2184), .A1N(n2134), 
        .Y(n3162) );
  AOI2BB2XL U2417 ( .B0(EX_data1[10]), .B1(n2137), .A0N(n2202), .A1N(n2134), 
        .Y(n3180) );
  AOI2BB2XL U2418 ( .B0(EX_data1[3]), .B1(n2137), .A0N(n2154), .A1N(n2134), 
        .Y(n3132) );
  AOI2BB2XL U2419 ( .B0(EX_data1[21]), .B1(n2137), .A0N(n2178), .A1N(n2134), 
        .Y(n3156) );
  AOI2BB2XL U2420 ( .B0(EX_data1[13]), .B1(n2137), .A0N(n2196), .A1N(n2134), 
        .Y(n3174) );
  AOI2BB2XL U2421 ( .B0(EX_data1[11]), .B1(n2137), .A0N(n2200), .A1N(n2134), 
        .Y(n3178) );
  AOI2BB2XL U2422 ( .B0(EX_data1[20]), .B1(n2137), .A0N(n2180), .A1N(n2134), 
        .Y(n3158) );
  AOI2BB2XL U2423 ( .B0(EX_data1[12]), .B1(n2137), .A0N(n2198), .A1N(n2134), 
        .Y(n3176) );
  AOI2BB2XL U2424 ( .B0(EX_data1[22]), .B1(n2137), .A0N(n2176), .A1N(n2134), 
        .Y(n3154) );
  AOI2BB2XL U2425 ( .B0(EX_data1[8]), .B1(n2137), .A0N(n2144), .A1N(n2134), 
        .Y(n3122) );
  AOI2BB2XL U2426 ( .B0(EX_data1[18]), .B1(n2137), .A0N(n2186), .A1N(n2134), 
        .Y(n3164) );
  AOI2BB2XL U2427 ( .B0(EX_data1[14]), .B1(n2137), .A0N(n2194), .A1N(n2134), 
        .Y(n3172) );
  AOI2BB2XL U2428 ( .B0(EX_data1[28]), .B1(n2137), .A0N(n2164), .A1N(n2134), 
        .Y(n3142) );
  AOI2BB2XL U2429 ( .B0(EX_data1[2]), .B1(n2137), .A0N(n2160), .A1N(n2134), 
        .Y(n3138) );
  AOI2BB2XL U2430 ( .B0(EX_data1[29]), .B1(n2137), .A0N(n2162), .A1N(n2134), 
        .Y(n3140) );
  AOI2BB2XL U2431 ( .B0(EX_data1[23]), .B1(n2137), .A0N(n2174), .A1N(n2134), 
        .Y(n3152) );
  AOI2BB2XL U2432 ( .B0(EX_data1[5]), .B1(n2137), .A0N(n2150), .A1N(n2134), 
        .Y(n3128) );
  AOI2BB2XL U2433 ( .B0(EX_data1[15]), .B1(n2137), .A0N(n2192), .A1N(n2134), 
        .Y(n3170) );
  AOI2BB2XL U2434 ( .B0(EX_data1[1]), .B1(n2137), .A0N(n2182), .A1N(n2134), 
        .Y(n3160) );
  AOI2BB2XL U2435 ( .B0(EX_data1[24]), .B1(n2137), .A0N(n2172), .A1N(n2134), 
        .Y(n3150) );
  AOI2BB2XL U2436 ( .B0(EX_data1[25]), .B1(n2137), .A0N(n2170), .A1N(n2134), 
        .Y(n3148) );
  AOI2BB2XL U2437 ( .B0(EX_data1[4]), .B1(n2137), .A0N(n2152), .A1N(n2134), 
        .Y(n3130) );
  AOI2BB2XL U2438 ( .B0(EX_data1[6]), .B1(n2137), .A0N(n2148), .A1N(n2134), 
        .Y(n3126) );
  AOI2BB2XL U2439 ( .B0(EX_data1[7]), .B1(n2137), .A0N(n2146), .A1N(n2134), 
        .Y(n3124) );
  AOI2BB2XL U2440 ( .B0(EX_data1[16]), .B1(n2137), .A0N(n2190), .A1N(n2134), 
        .Y(n3168) );
  AOI2BB2XL U2441 ( .B0(EX_data1[17]), .B1(n2137), .A0N(n2188), .A1N(n2134), 
        .Y(n3166) );
  AOI2BB2XL U2442 ( .B0(EX_data1[0]), .B1(n2137), .A0N(n2204), .A1N(n2134), 
        .Y(n3182) );
  AOI2BB2XL U2443 ( .B0(EX_data1[30]), .B1(n2137), .A0N(n2158), .A1N(n2134), 
        .Y(n3136) );
  AOI2BB2XL U2444 ( .B0(EX_data1[31]), .B1(n2137), .A0N(n2156), .A1N(n2134), 
        .Y(n3134) );
  NAND2XL U2445 ( .A(BranchAddr[6]), .B(n3036), .Y(n3047) );
  OAI211XL U2446 ( .A0(n3248), .A1(n2139), .B0(n3041), .C0(n3042), .Y(n1351)
         );
  NAND2XL U2447 ( .A(BranchAddr[3]), .B(n3036), .Y(n3041) );
  OAI211XL U2448 ( .A0(n3221), .A1(n2139), .B0(n3095), .C0(n3096), .Y(n1324)
         );
  NAND2XL U2449 ( .A(BranchAddr[30]), .B(n3036), .Y(n3095) );
  OAI211XL U2450 ( .A0(n3222), .A1(n2139), .B0(n3093), .C0(n3094), .Y(n1325)
         );
  NAND2XL U2451 ( .A(BranchAddr[29]), .B(n3036), .Y(n3093) );
  OAI211XL U2452 ( .A0(n3223), .A1(n2139), .B0(n3091), .C0(n3092), .Y(n1326)
         );
  NAND2XL U2453 ( .A(BranchAddr[28]), .B(n3036), .Y(n3091) );
  OAI211XL U2454 ( .A0(n3224), .A1(n2139), .B0(n3089), .C0(n3090), .Y(n1327)
         );
  NAND2XL U2455 ( .A(BranchAddr[27]), .B(n3036), .Y(n3089) );
  OAI211XL U2456 ( .A0(n3225), .A1(n2139), .B0(n3087), .C0(n3088), .Y(n1328)
         );
  NAND2XL U2457 ( .A(BranchAddr[26]), .B(n3036), .Y(n3087) );
  OAI211XL U2458 ( .A0(n3226), .A1(n2139), .B0(n3085), .C0(n3086), .Y(n1329)
         );
  NAND2XL U2459 ( .A(BranchAddr[25]), .B(n3036), .Y(n3085) );
  OAI211XL U2460 ( .A0(n3227), .A1(n2139), .B0(n3083), .C0(n3084), .Y(n1330)
         );
  NAND2XL U2461 ( .A(BranchAddr[24]), .B(n3036), .Y(n3083) );
  OAI211XL U2462 ( .A0(n3228), .A1(n2139), .B0(n3081), .C0(n3082), .Y(n1331)
         );
  NAND2XL U2463 ( .A(BranchAddr[23]), .B(n3036), .Y(n3081) );
  OAI211XL U2464 ( .A0(n3229), .A1(n2139), .B0(n3079), .C0(n3080), .Y(n1332)
         );
  NAND2XL U2465 ( .A(BranchAddr[22]), .B(n3036), .Y(n3079) );
  OAI211XL U2466 ( .A0(n3230), .A1(n2139), .B0(n3077), .C0(n3078), .Y(n1333)
         );
  NAND2XL U2467 ( .A(BranchAddr[21]), .B(n3036), .Y(n3077) );
  OAI211XL U2468 ( .A0(n3231), .A1(n2139), .B0(n3075), .C0(n3076), .Y(n1334)
         );
  NAND2XL U2469 ( .A(BranchAddr[20]), .B(n3036), .Y(n3075) );
  OAI211XL U2470 ( .A0(n3232), .A1(n2139), .B0(n3073), .C0(n3074), .Y(n1335)
         );
  NAND2XL U2471 ( .A(BranchAddr[19]), .B(n3036), .Y(n3073) );
  OAI211XL U2472 ( .A0(n3233), .A1(n2139), .B0(n3071), .C0(n3072), .Y(n1336)
         );
  NAND2XL U2473 ( .A(BranchAddr[18]), .B(n3036), .Y(n3071) );
  OAI211XL U2474 ( .A0(n3234), .A1(n2139), .B0(n3069), .C0(n3070), .Y(n1337)
         );
  NAND2XL U2475 ( .A(BranchAddr[17]), .B(n3036), .Y(n3069) );
  OAI211XL U2476 ( .A0(n3235), .A1(n2139), .B0(n3067), .C0(n3068), .Y(n1338)
         );
  NAND2XL U2477 ( .A(BranchAddr[16]), .B(n3036), .Y(n3067) );
  OAI211XL U2478 ( .A0(n3236), .A1(n2139), .B0(n3065), .C0(n3066), .Y(n1339)
         );
  NAND2XL U2479 ( .A(BranchAddr[15]), .B(n3036), .Y(n3065) );
  OAI211XL U2480 ( .A0(n3237), .A1(n2139), .B0(n3063), .C0(n3064), .Y(n1340)
         );
  NAND2XL U2481 ( .A(BranchAddr[14]), .B(n3036), .Y(n3063) );
  OAI211XL U2482 ( .A0(n3238), .A1(n2139), .B0(n3061), .C0(n3062), .Y(n1341)
         );
  NAND2XL U2483 ( .A(BranchAddr[13]), .B(n3036), .Y(n3061) );
  OAI211XL U2484 ( .A0(n3239), .A1(n2139), .B0(n3059), .C0(n3060), .Y(n1342)
         );
  NAND2XL U2485 ( .A(BranchAddr[12]), .B(n3036), .Y(n3059) );
  OAI211XL U2486 ( .A0(n3240), .A1(n2139), .B0(n3057), .C0(n3058), .Y(n1343)
         );
  NAND2XL U2487 ( .A(BranchAddr[11]), .B(n3036), .Y(n3057) );
  OAI211XL U2488 ( .A0(n3241), .A1(n2139), .B0(n3055), .C0(n3056), .Y(n1344)
         );
  NAND2XL U2489 ( .A(BranchAddr[10]), .B(n3036), .Y(n3055) );
  OAI211XL U2490 ( .A0(n3242), .A1(n2139), .B0(n3053), .C0(n3054), .Y(n1345)
         );
  NAND2XL U2491 ( .A(BranchAddr[9]), .B(n3036), .Y(n3053) );
  OAI211XL U2492 ( .A0(n3243), .A1(n2139), .B0(n3051), .C0(n3052), .Y(n1346)
         );
  NAND2XL U2493 ( .A(BranchAddr[8]), .B(n3036), .Y(n3051) );
  OAI211XL U2494 ( .A0(n3244), .A1(n2139), .B0(n3049), .C0(n3050), .Y(n1347)
         );
  NAND2XL U2495 ( .A(BranchAddr[7]), .B(n3036), .Y(n3049) );
  OAI211XL U2496 ( .A0(n3246), .A1(n2139), .B0(n3045), .C0(n3046), .Y(n1349)
         );
  NAND2XL U2497 ( .A(BranchAddr[5]), .B(n3036), .Y(n3045) );
  OAI211XL U2498 ( .A0(n3247), .A1(n2139), .B0(n3043), .C0(n3044), .Y(n1350)
         );
  NAND2XL U2499 ( .A(BranchAddr[4]), .B(n3036), .Y(n3043) );
  OAI211XL U2500 ( .A0(n3250), .A1(n2139), .B0(n3037), .C0(n3038), .Y(n1353)
         );
  NAND2XL U2501 ( .A(BranchAddr[1]), .B(n3036), .Y(n3037) );
  AOI22XL U2502 ( .A0(PC_plus4[1]), .A1(n3035), .B0(read_data1[1]), .B1(n2132), 
        .Y(n3038) );
  OAI211XL U2503 ( .A0(n3251), .A1(n2139), .B0(n3033), .C0(n3034), .Y(n1354)
         );
  NAND2XL U2504 ( .A(BranchAddr[0]), .B(n3036), .Y(n3033) );
  AOI22XL U2505 ( .A0(PC_plus4[0]), .A1(n3035), .B0(read_data1[0]), .B1(n2132), 
        .Y(n3034) );
  AND3X2 U2506 ( .A(WB_WB[0]), .B(WB_Rd[3]), .C(WB_Rd[4]), .Y(n3103) );
  AND3X2 U2507 ( .A(WB_WB[0]), .B(n3015), .C(WB_Rd[4]), .Y(n2993) );
  AOI2BB2XL U2508 ( .B0(EX_data2[15]), .B1(n2138), .A0N(n2192), .A1N(n2206), 
        .Y(n3213) );
  AOI2BB2XL U2509 ( .B0(EX_data2[16]), .B1(n2138), .A0N(n2190), .A1N(n2206), 
        .Y(n3212) );
  AOI2BB2XL U2510 ( .B0(EX_data2[3]), .B1(n2138), .A0N(n2154), .A1N(n2206), 
        .Y(n3194) );
  AOI2BB2XL U2511 ( .B0(EX_data2[5]), .B1(n2138), .A0N(n2150), .A1N(n2206), 
        .Y(n3192) );
  AOI2BB2XL U2512 ( .B0(EX_data2[4]), .B1(n2138), .A0N(n2152), .A1N(n2206), 
        .Y(n3193) );
  AOI2BB2XL U2513 ( .B0(EX_data2[1]), .B1(n2138), .A0N(n2182), .A1N(n2206), 
        .Y(n3208) );
  AOI2BB2XL U2514 ( .B0(EX_data2[0]), .B1(n2138), .A0N(n2204), .A1N(n2206), 
        .Y(n3219) );
  AOI2BB2XL U2515 ( .B0(EX_data2[2]), .B1(n2138), .A0N(n2160), .A1N(n2206), 
        .Y(n3197) );
  AOI2BB2XL U2516 ( .B0(EX_data2[10]), .B1(n2138), .A0N(n2202), .A1N(n2206), 
        .Y(n3218) );
  AOI2BB2XL U2517 ( .B0(EX_data2[11]), .B1(n2138), .A0N(n2200), .A1N(n2206), 
        .Y(n3217) );
  AOI2BB2XL U2518 ( .B0(EX_data2[13]), .B1(n2138), .A0N(n2196), .A1N(n2206), 
        .Y(n3215) );
  AOI2BB2XL U2519 ( .B0(EX_data2[8]), .B1(n2138), .A0N(n2144), .A1N(n2206), 
        .Y(n3189) );
  AOI2BB2XL U2520 ( .B0(EX_data2[14]), .B1(n2138), .A0N(n2194), .A1N(n2206), 
        .Y(n3214) );
  AOI2BB2XL U2521 ( .B0(EX_data2[25]), .B1(n2138), .A0N(n2170), .A1N(n2206), 
        .Y(n3202) );
  AOI2BB2XL U2522 ( .B0(EX_data2[6]), .B1(n2138), .A0N(n2148), .A1N(n2206), 
        .Y(n3191) );
  AOI2BB2XL U2523 ( .B0(EX_data2[7]), .B1(n2138), .A0N(n2146), .A1N(n2206), 
        .Y(n3190) );
  AOI2BB2XL U2524 ( .B0(EX_data2[12]), .B1(n2138), .A0N(n2198), .A1N(n2206), 
        .Y(n3216) );
  AOI2BB2XL U2525 ( .B0(EX_data2[31]), .B1(n2138), .A0N(n2156), .A1N(n2206), 
        .Y(n3195) );
  AOI2BB2XL U2526 ( .B0(EX_data2[18]), .B1(n2138), .A0N(n2186), .A1N(n2206), 
        .Y(n3210) );
  AOI2BB2XL U2527 ( .B0(EX_data2[30]), .B1(n2138), .A0N(n2158), .A1N(n2206), 
        .Y(n3196) );
  AOI2BB2XL U2528 ( .B0(EX_data2[9]), .B1(n2138), .A0N(n2142), .A1N(n2206), 
        .Y(n3184) );
  AOI2BB2XL U2529 ( .B0(EX_data2[26]), .B1(n2138), .A0N(n2168), .A1N(n2206), 
        .Y(n3201) );
  AOI2BB2XL U2530 ( .B0(EX_data2[27]), .B1(n2138), .A0N(n2166), .A1N(n2206), 
        .Y(n3200) );
  AOI2BB2XL U2531 ( .B0(EX_data2[28]), .B1(n2138), .A0N(n2164), .A1N(n2206), 
        .Y(n3199) );
  AOI2BB2XL U2532 ( .B0(EX_data2[17]), .B1(n2138), .A0N(n2188), .A1N(n2206), 
        .Y(n3211) );
  AOI2BB2XL U2533 ( .B0(EX_data2[29]), .B1(n2138), .A0N(n2162), .A1N(n2206), 
        .Y(n3198) );
  AOI2BB2XL U2534 ( .B0(EX_data2[24]), .B1(n2138), .A0N(n2172), .A1N(n2206), 
        .Y(n3203) );
  AOI2BB2XL U2535 ( .B0(EX_data2[22]), .B1(n2138), .A0N(n2176), .A1N(n2206), 
        .Y(n3205) );
  AOI2BB2XL U2536 ( .B0(EX_data2[23]), .B1(n2138), .A0N(n2174), .A1N(n2206), 
        .Y(n3204) );
  AOI2BB2XL U2537 ( .B0(EX_data2[19]), .B1(n2138), .A0N(n2184), .A1N(n2206), 
        .Y(n3209) );
  AOI2BB2XL U2538 ( .B0(EX_data2[20]), .B1(n2138), .A0N(n2180), .A1N(n2206), 
        .Y(n3207) );
  AOI2BB2XL U2539 ( .B0(EX_data2[21]), .B1(n2138), .A0N(n2178), .A1N(n2206), 
        .Y(n3206) );
  MXI2XL U2540 ( .A(n2619), .B(n2620), .S0(N77), .Y(read_data2[6]) );
  MXI2XL U2541 ( .A(n2663), .B(n2664), .S0(N77), .Y(read_data2[28]) );
  MXI2XL U2542 ( .A(n2665), .B(n2666), .S0(N77), .Y(read_data2[29]) );
  MXI2XL U2543 ( .A(n2667), .B(n2668), .S0(N77), .Y(read_data2[30]) );
  MXI2XL U2544 ( .A(n2669), .B(n2670), .S0(N77), .Y(read_data2[31]) );
  MXI2XL U2545 ( .A(n2621), .B(n2622), .S0(N77), .Y(read_data2[7]) );
  MXI2XL U2546 ( .A(n2623), .B(n2624), .S0(N77), .Y(read_data2[8]) );
  MXI2XL U2547 ( .A(n2625), .B(n2626), .S0(N77), .Y(read_data2[9]) );
  MXI2XL U2548 ( .A(n2627), .B(n2628), .S0(N77), .Y(read_data2[10]) );
  MXI2XL U2549 ( .A(n2629), .B(n2630), .S0(N77), .Y(read_data2[11]) );
  MXI2XL U2550 ( .A(n2631), .B(n2632), .S0(N77), .Y(read_data2[12]) );
  MXI2XL U2551 ( .A(n2633), .B(n2634), .S0(N77), .Y(read_data2[13]) );
  MXI2XL U2552 ( .A(n2635), .B(n2636), .S0(N77), .Y(read_data2[14]) );
  MXI2XL U2553 ( .A(n2637), .B(n2638), .S0(N77), .Y(read_data2[15]) );
  MXI2XL U2554 ( .A(n2639), .B(n2640), .S0(N77), .Y(read_data2[16]) );
  MXI2XL U2555 ( .A(n2641), .B(n2642), .S0(N77), .Y(read_data2[17]) );
  MXI2XL U2556 ( .A(n2643), .B(n2644), .S0(N77), .Y(read_data2[18]) );
  MXI2XL U2557 ( .A(n2645), .B(n2646), .S0(N77), .Y(read_data2[19]) );
  MXI2XL U2558 ( .A(n2647), .B(n2648), .S0(N77), .Y(read_data2[20]) );
  MXI2XL U2559 ( .A(n2649), .B(n2650), .S0(N77), .Y(read_data2[21]) );
  MXI2XL U2560 ( .A(n2651), .B(n2652), .S0(N77), .Y(read_data2[22]) );
  MXI2XL U2561 ( .A(n2653), .B(n2654), .S0(N77), .Y(read_data2[23]) );
  MXI2XL U2562 ( .A(n2655), .B(n2656), .S0(N77), .Y(read_data2[24]) );
  MXI2XL U2563 ( .A(n2657), .B(n2658), .S0(N77), .Y(read_data2[25]) );
  MXI2XL U2564 ( .A(n2659), .B(n2660), .S0(N77), .Y(read_data2[26]) );
  MXI2XL U2565 ( .A(n2661), .B(n2662), .S0(N77), .Y(read_data2[27]) );
  MX2X1 U2566 ( .A(after_B_mux[11]), .B(EX_signextend[11]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[11]) );
  MX2X1 U2567 ( .A(after_B_mux[13]), .B(EX_signextend[13]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[13]) );
  MX2X1 U2568 ( .A(after_B_mux[9]), .B(EX_signextend[9]), .S0(EX_reg[3]), .Y(
        after_ALUSrc[9]) );
  MX2X1 U2569 ( .A(after_B_mux[27]), .B(EX_signextend[27]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[27]) );
  MX2X1 U2570 ( .A(after_B_mux[10]), .B(EX_signextend[10]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[10]) );
  MX2X1 U2571 ( .A(after_B_mux[26]), .B(EX_signextend[26]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[26]) );
  MX2X1 U2572 ( .A(after_B_mux[28]), .B(EX_signextend[28]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[28]) );
  MX2X1 U2573 ( .A(after_B_mux[12]), .B(EX_signextend[12]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[12]) );
  MX2X1 U2574 ( .A(after_B_mux[20]), .B(EX_signextend[20]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[20]) );
  MX2X1 U2575 ( .A(after_B_mux[19]), .B(EX_signextend[19]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[19]) );
  MX2X1 U2576 ( .A(after_B_mux[21]), .B(EX_signextend[21]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[21]) );
  MX2X1 U2577 ( .A(after_B_mux[29]), .B(EX_signextend[29]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[29]) );
  NOR2BXL U2578 ( .AN(ALUOp[1]), .B(n3116), .Y(EX_after_detect[1]) );
  NOR2BXL U2579 ( .AN(ALUOp[0]), .B(n3116), .Y(EX_after_detect[0]) );
  NOR2BXL U2580 ( .AN(M[2]), .B(n3116), .Y(MEM_after_detect[2]) );
  NOR2BXL U2581 ( .AN(\WB[0] ), .B(n3116), .Y(WB_after_detect[0]) );
  CLKBUFX3 U2582 ( .A(n70), .Y(n2209) );
  CLKBUFX3 U2583 ( .A(N74), .Y(n2222) );
  BUFX12 U2584 ( .A(n2286), .Y(n2283) );
  BUFX12 U2585 ( .A(n2286), .Y(n2282) );
  BUFX12 U2586 ( .A(n2286), .Y(n2278) );
  BUFX12 U2587 ( .A(n2286), .Y(n2284) );
  BUFX12 U2588 ( .A(n2286), .Y(n2271) );
  BUFX12 U2589 ( .A(n2286), .Y(n2272) );
  BUFX12 U2590 ( .A(n2286), .Y(n2273) );
  BUFX12 U2591 ( .A(n2286), .Y(n2274) );
  BUFX12 U2592 ( .A(rst_n), .Y(n2275) );
  BUFX12 U2593 ( .A(n2286), .Y(n2276) );
  BUFX12 U2594 ( .A(n2286), .Y(n2277) );
  BUFX12 U2595 ( .A(n2285), .Y(n2279) );
  BUFX12 U2596 ( .A(rst_n), .Y(n2280) );
  BUFX12 U2597 ( .A(n2286), .Y(n2281) );
  CLKBUFX8 U2598 ( .A(n2286), .Y(n2285) );
  BUFX4 U2599 ( .A(N69), .Y(n2247) );
  BUFX4 U2600 ( .A(n2252), .Y(n2248) );
  BUFX4 U2601 ( .A(N69), .Y(n2249) );
  BUFX4 U2602 ( .A(n2242), .Y(n2250) );
  BUFX4 U2603 ( .A(n2252), .Y(n2243) );
  BUFX4 U2604 ( .A(N69), .Y(n2244) );
  BUFX4 U2605 ( .A(N69), .Y(n2245) );
  BUFX4 U2606 ( .A(N69), .Y(n2246) );
  CLKBUFX3 U2607 ( .A(n2233), .Y(n2234) );
  CLKBUFX3 U2608 ( .A(n2227), .Y(n2235) );
  CLKBUFX3 U2609 ( .A(n2233), .Y(n2236) );
  CLKBUFX3 U2610 ( .A(n2232), .Y(n2237) );
  CLKBUFX3 U2611 ( .A(N73), .Y(n2238) );
  CLKBUFX3 U2612 ( .A(n2240), .Y(n2239) );
  CLKBUFX3 U2613 ( .A(n2238), .Y(n2240) );
  CLKBUFX3 U2614 ( .A(n2228), .Y(n2241) );
  CLKBUFX3 U2615 ( .A(N73), .Y(n2225) );
  CLKBUFX3 U2616 ( .A(n2227), .Y(n2226) );
  CLKBUFX3 U2617 ( .A(N73), .Y(n2227) );
  CLKBUFX3 U2618 ( .A(n2238), .Y(n2228) );
  CLKBUFX3 U2619 ( .A(n2233), .Y(n2229) );
  CLKBUFX3 U2620 ( .A(N73), .Y(n2230) );
  CLKBUFX3 U2621 ( .A(n2225), .Y(n2231) );
  CLKBUFX3 U2622 ( .A(N73), .Y(n2233) );
  CLKBUFX3 U2623 ( .A(N73), .Y(n2232) );
  CLKBUFX3 U2624 ( .A(n2254), .Y(n2263) );
  CLKBUFX3 U2625 ( .A(n2262), .Y(n2264) );
  CLKBUFX3 U2626 ( .A(n2254), .Y(n2265) );
  CLKBUFX3 U2627 ( .A(n2256), .Y(n2266) );
  CLKBUFX3 U2628 ( .A(n2253), .Y(n2267) );
  CLKBUFX3 U2629 ( .A(n2255), .Y(n2268) );
  CLKBUFX3 U2630 ( .A(n2261), .Y(n2269) );
  CLKBUFX3 U2631 ( .A(n2266), .Y(n2270) );
  CLKBUFX3 U2632 ( .A(N68), .Y(n2254) );
  CLKBUFX3 U2633 ( .A(n2256), .Y(n2255) );
  CLKBUFX3 U2634 ( .A(N68), .Y(n2256) );
  CLKBUFX3 U2635 ( .A(n2261), .Y(n2257) );
  CLKBUFX3 U2636 ( .A(n2253), .Y(n2258) );
  CLKBUFX3 U2637 ( .A(N68), .Y(n2259) );
  CLKBUFX3 U2638 ( .A(n2253), .Y(n2260) );
  CLKBUFX3 U2639 ( .A(N68), .Y(n2262) );
  CLKBUFX3 U2640 ( .A(N68), .Y(n2261) );
  CLKBUFX3 U2641 ( .A(n2223), .Y(n2217) );
  CLKBUFX3 U2642 ( .A(n2223), .Y(n2218) );
  CLKBUFX3 U2643 ( .A(n2223), .Y(n2219) );
  CLKBUFX3 U2644 ( .A(N74), .Y(n2220) );
  CLKBUFX3 U2645 ( .A(N74), .Y(n2221) );
  CLKBUFX3 U2646 ( .A(n2223), .Y(n2211) );
  CLKBUFX3 U2647 ( .A(n2223), .Y(n2212) );
  CLKBUFX3 U2648 ( .A(n2223), .Y(n2213) );
  CLKBUFX3 U2649 ( .A(n2223), .Y(n2214) );
  CLKBUFX3 U2650 ( .A(N74), .Y(n2215) );
  CLKBUFX3 U2651 ( .A(n2223), .Y(n2216) );
  CLKBUFX3 U2652 ( .A(n2223), .Y(n2210) );
  MXI4XL U2653 ( .A(\reg_file_next[4][0] ), .B(\reg_file_next[5][0] ), .C(
        \reg_file_next[6][0] ), .D(\reg_file_next[7][0] ), .S0(n2233), .S1(
        n2216), .Y(n2677) );
  MXI4XL U2654 ( .A(\reg_file_next[20][0] ), .B(\reg_file_next[21][0] ), .C(
        \reg_file_next[22][0] ), .D(\reg_file_next[23][0] ), .S0(n2233), .S1(
        n2216), .Y(n2673) );
  MXI4XL U2655 ( .A(\reg_file_next[4][1] ), .B(\reg_file_next[5][1] ), .C(
        \reg_file_next[6][1] ), .D(\reg_file_next[7][1] ), .S0(n2234), .S1(
        n2217), .Y(n2685) );
  MXI4XL U2656 ( .A(\reg_file_next[20][1] ), .B(\reg_file_next[21][1] ), .C(
        \reg_file_next[22][1] ), .D(\reg_file_next[23][1] ), .S0(n2234), .S1(
        n2217), .Y(n2681) );
  MXI4XL U2657 ( .A(\reg_file_next[4][2] ), .B(\reg_file_next[5][2] ), .C(
        \reg_file_next[6][2] ), .D(\reg_file_next[7][2] ), .S0(n2234), .S1(
        n2217), .Y(n2693) );
  MXI4XL U2658 ( .A(\reg_file_next[20][2] ), .B(\reg_file_next[21][2] ), .C(
        \reg_file_next[22][2] ), .D(\reg_file_next[23][2] ), .S0(n2234), .S1(
        n2217), .Y(n2689) );
  MXI4XL U2659 ( .A(\reg_file_next[4][3] ), .B(\reg_file_next[5][3] ), .C(
        \reg_file_next[6][3] ), .D(\reg_file_next[7][3] ), .S0(n2235), .S1(
        n2218), .Y(n2701) );
  MXI4XL U2660 ( .A(\reg_file_next[20][3] ), .B(\reg_file_next[21][3] ), .C(
        \reg_file_next[22][3] ), .D(\reg_file_next[23][3] ), .S0(n2235), .S1(
        n2217), .Y(n2697) );
  MXI4XL U2661 ( .A(\reg_file_next[4][4] ), .B(\reg_file_next[5][4] ), .C(
        \reg_file_next[6][4] ), .D(\reg_file_next[7][4] ), .S0(n2236), .S1(
        n2218), .Y(n2709) );
  MXI4XL U2662 ( .A(\reg_file_next[20][4] ), .B(\reg_file_next[21][4] ), .C(
        \reg_file_next[22][4] ), .D(\reg_file_next[23][4] ), .S0(n2235), .S1(
        n2218), .Y(n2705) );
  MXI4XL U2663 ( .A(\reg_file_next[4][5] ), .B(\reg_file_next[5][5] ), .C(
        \reg_file_next[6][5] ), .D(\reg_file_next[7][5] ), .S0(n2236), .S1(
        n2218), .Y(n2717) );
  MXI4XL U2664 ( .A(\reg_file_next[20][5] ), .B(\reg_file_next[21][5] ), .C(
        \reg_file_next[22][5] ), .D(\reg_file_next[23][5] ), .S0(n2236), .S1(
        n2218), .Y(n2713) );
  MXI4XL U2665 ( .A(\reg_file_next[4][6] ), .B(\reg_file_next[5][6] ), .C(
        \reg_file_next[6][6] ), .D(\reg_file_next[7][6] ), .S0(n2237), .S1(
        n2219), .Y(n2725) );
  MXI4XL U2666 ( .A(\reg_file_next[20][6] ), .B(\reg_file_next[21][6] ), .C(
        \reg_file_next[22][6] ), .D(\reg_file_next[23][6] ), .S0(n2236), .S1(
        n2219), .Y(n2721) );
  MXI4XL U2667 ( .A(\reg_file_next[4][7] ), .B(\reg_file_next[5][7] ), .C(
        \reg_file_next[6][7] ), .D(\reg_file_next[7][7] ), .S0(n2237), .S1(
        n2219), .Y(n2733) );
  MXI4XL U2668 ( .A(\reg_file_next[20][7] ), .B(\reg_file_next[21][7] ), .C(
        \reg_file_next[22][7] ), .D(\reg_file_next[23][7] ), .S0(n2237), .S1(
        n2219), .Y(n2729) );
  MXI4XL U2669 ( .A(\reg_file_next[4][8] ), .B(\reg_file_next[5][8] ), .C(
        \reg_file_next[6][8] ), .D(\reg_file_next[7][8] ), .S0(n2238), .S1(
        n2220), .Y(n2741) );
  MXI4XL U2670 ( .A(\reg_file_next[20][8] ), .B(\reg_file_next[21][8] ), .C(
        \reg_file_next[22][8] ), .D(\reg_file_next[23][8] ), .S0(n2238), .S1(
        n2220), .Y(n2737) );
  MXI4XL U2671 ( .A(\reg_file_next[4][9] ), .B(\reg_file_next[5][9] ), .C(
        \reg_file_next[6][9] ), .D(\reg_file_next[7][9] ), .S0(n2239), .S1(
        n2220), .Y(n2749) );
  MXI4XL U2672 ( .A(\reg_file_next[20][9] ), .B(\reg_file_next[21][9] ), .C(
        \reg_file_next[22][9] ), .D(\reg_file_next[23][9] ), .S0(n2238), .S1(
        n2220), .Y(n2745) );
  MXI4XL U2673 ( .A(\reg_file_next[4][10] ), .B(\reg_file_next[5][10] ), .C(
        \reg_file_next[6][10] ), .D(\reg_file_next[7][10] ), .S0(n2239), .S1(
        n2221), .Y(n2757) );
  MXI4XL U2674 ( .A(\reg_file_next[20][10] ), .B(\reg_file_next[21][10] ), .C(
        \reg_file_next[22][10] ), .D(\reg_file_next[23][10] ), .S0(n2239), 
        .S1(n2220), .Y(n2753) );
  MXI4XL U2675 ( .A(\reg_file_next[4][11] ), .B(\reg_file_next[5][11] ), .C(
        \reg_file_next[6][11] ), .D(\reg_file_next[7][11] ), .S0(n2240), .S1(
        n2221), .Y(n2765) );
  MXI4XL U2676 ( .A(\reg_file_next[20][11] ), .B(\reg_file_next[21][11] ), .C(
        \reg_file_next[22][11] ), .D(\reg_file_next[23][11] ), .S0(n2239), 
        .S1(n2221), .Y(n2761) );
  MXI4XL U2677 ( .A(\reg_file_next[4][12] ), .B(\reg_file_next[5][12] ), .C(
        \reg_file_next[6][12] ), .D(\reg_file_next[7][12] ), .S0(n2240), .S1(
        n2221), .Y(n2773) );
  MXI4XL U2678 ( .A(\reg_file_next[20][12] ), .B(\reg_file_next[21][12] ), .C(
        \reg_file_next[22][12] ), .D(\reg_file_next[23][12] ), .S0(n2240), 
        .S1(n2221), .Y(n2769) );
  MXI4XL U2679 ( .A(\reg_file_next[4][13] ), .B(\reg_file_next[5][13] ), .C(
        \reg_file_next[6][13] ), .D(\reg_file_next[7][13] ), .S0(n2241), .S1(
        n2222), .Y(n2781) );
  MXI4XL U2680 ( .A(\reg_file_next[20][13] ), .B(\reg_file_next[21][13] ), .C(
        \reg_file_next[22][13] ), .D(\reg_file_next[23][13] ), .S0(n2241), 
        .S1(n2222), .Y(n2777) );
  MXI4XL U2681 ( .A(\reg_file_next[4][14] ), .B(\reg_file_next[5][14] ), .C(
        \reg_file_next[6][14] ), .D(\reg_file_next[7][14] ), .S0(n2241), .S1(
        n2222), .Y(n2789) );
  MXI4XL U2682 ( .A(\reg_file_next[20][14] ), .B(\reg_file_next[21][14] ), .C(
        \reg_file_next[22][14] ), .D(\reg_file_next[23][14] ), .S0(n2241), 
        .S1(n2222), .Y(n2785) );
  MXI4XL U2683 ( .A(\reg_file_next[4][15] ), .B(\reg_file_next[5][15] ), .C(
        \reg_file_next[6][15] ), .D(\reg_file_next[7][15] ), .S0(n2234), .S1(
        N74), .Y(n2797) );
  MXI4XL U2684 ( .A(\reg_file_next[20][15] ), .B(\reg_file_next[21][15] ), .C(
        \reg_file_next[22][15] ), .D(\reg_file_next[23][15] ), .S0(n2235), 
        .S1(n2222), .Y(n2793) );
  MXI4XL U2685 ( .A(\reg_file_next[4][16] ), .B(\reg_file_next[5][16] ), .C(
        \reg_file_next[6][16] ), .D(\reg_file_next[7][16] ), .S0(n2224), .S1(
        n2210), .Y(n2805) );
  MXI4XL U2686 ( .A(\reg_file_next[20][16] ), .B(\reg_file_next[21][16] ), .C(
        \reg_file_next[22][16] ), .D(\reg_file_next[23][16] ), .S0(n2224), 
        .S1(n2210), .Y(n2801) );
  MXI4XL U2687 ( .A(\reg_file_next[4][17] ), .B(\reg_file_next[5][17] ), .C(
        \reg_file_next[6][17] ), .D(\reg_file_next[7][17] ), .S0(n2225), .S1(
        n2211), .Y(n2813) );
  MXI4XL U2688 ( .A(\reg_file_next[20][17] ), .B(\reg_file_next[21][17] ), .C(
        \reg_file_next[22][17] ), .D(\reg_file_next[23][17] ), .S0(n2225), 
        .S1(n2210), .Y(n2809) );
  MXI4XL U2689 ( .A(\reg_file_next[4][18] ), .B(\reg_file_next[5][18] ), .C(
        \reg_file_next[6][18] ), .D(\reg_file_next[7][18] ), .S0(n2225), .S1(
        n2211), .Y(n2821) );
  MXI4XL U2690 ( .A(\reg_file_next[20][18] ), .B(\reg_file_next[21][18] ), .C(
        \reg_file_next[22][18] ), .D(\reg_file_next[23][18] ), .S0(n2225), 
        .S1(n2211), .Y(n2817) );
  MXI4XL U2691 ( .A(\reg_file_next[4][19] ), .B(\reg_file_next[5][19] ), .C(
        \reg_file_next[6][19] ), .D(\reg_file_next[7][19] ), .S0(n2226), .S1(
        n2211), .Y(n2829) );
  MXI4XL U2692 ( .A(\reg_file_next[20][19] ), .B(\reg_file_next[21][19] ), .C(
        \reg_file_next[22][19] ), .D(\reg_file_next[23][19] ), .S0(n2226), 
        .S1(n2211), .Y(n2825) );
  MXI4XL U2693 ( .A(\reg_file_next[4][20] ), .B(\reg_file_next[5][20] ), .C(
        \reg_file_next[6][20] ), .D(\reg_file_next[7][20] ), .S0(n2227), .S1(
        n2212), .Y(n2837) );
  MXI4XL U2694 ( .A(\reg_file_next[20][20] ), .B(\reg_file_next[21][20] ), .C(
        \reg_file_next[22][20] ), .D(\reg_file_next[23][20] ), .S0(n2226), 
        .S1(n2212), .Y(n2833) );
  MXI4XL U2695 ( .A(\reg_file_next[4][21] ), .B(\reg_file_next[5][21] ), .C(
        \reg_file_next[6][21] ), .D(\reg_file_next[7][21] ), .S0(n2227), .S1(
        n2212), .Y(n2845) );
  MXI4XL U2696 ( .A(\reg_file_next[20][21] ), .B(\reg_file_next[21][21] ), .C(
        \reg_file_next[22][21] ), .D(\reg_file_next[23][21] ), .S0(n2227), 
        .S1(n2212), .Y(n2841) );
  MXI4XL U2697 ( .A(\reg_file_next[4][22] ), .B(\reg_file_next[5][22] ), .C(
        \reg_file_next[6][22] ), .D(\reg_file_next[7][22] ), .S0(n2228), .S1(
        n2213), .Y(n2853) );
  MXI4XL U2698 ( .A(\reg_file_next[20][22] ), .B(\reg_file_next[21][22] ), .C(
        \reg_file_next[22][22] ), .D(\reg_file_next[23][22] ), .S0(n2227), 
        .S1(n2212), .Y(n2849) );
  MXI4XL U2699 ( .A(\reg_file_next[4][23] ), .B(\reg_file_next[5][23] ), .C(
        \reg_file_next[6][23] ), .D(\reg_file_next[7][23] ), .S0(n2228), .S1(
        n2213), .Y(n2861) );
  MXI4XL U2700 ( .A(\reg_file_next[20][23] ), .B(\reg_file_next[21][23] ), .C(
        \reg_file_next[22][23] ), .D(\reg_file_next[23][23] ), .S0(n2228), 
        .S1(n2213), .Y(n2857) );
  MXI4XL U2701 ( .A(\reg_file_next[4][24] ), .B(\reg_file_next[5][24] ), .C(
        \reg_file_next[6][24] ), .D(\reg_file_next[7][24] ), .S0(n2229), .S1(
        n2213), .Y(n2869) );
  MXI4XL U2702 ( .A(\reg_file_next[20][24] ), .B(\reg_file_next[21][24] ), .C(
        \reg_file_next[22][24] ), .D(\reg_file_next[23][24] ), .S0(n2229), 
        .S1(n2213), .Y(n2865) );
  MXI4XL U2703 ( .A(\reg_file_next[4][25] ), .B(\reg_file_next[5][25] ), .C(
        \reg_file_next[6][25] ), .D(\reg_file_next[7][25] ), .S0(n2229), .S1(
        n2214), .Y(n2877) );
  MXI4XL U2704 ( .A(\reg_file_next[20][25] ), .B(\reg_file_next[21][25] ), .C(
        \reg_file_next[22][25] ), .D(\reg_file_next[23][25] ), .S0(n2229), 
        .S1(n2214), .Y(n2873) );
  MXI4XL U2705 ( .A(\reg_file_next[4][26] ), .B(\reg_file_next[5][26] ), .C(
        \reg_file_next[6][26] ), .D(\reg_file_next[7][26] ), .S0(n2230), .S1(
        n2214), .Y(n2885) );
  MXI4XL U2706 ( .A(\reg_file_next[20][26] ), .B(\reg_file_next[21][26] ), .C(
        \reg_file_next[22][26] ), .D(\reg_file_next[23][26] ), .S0(n2230), 
        .S1(n2214), .Y(n2881) );
  MXI4XL U2707 ( .A(\reg_file_next[4][27] ), .B(\reg_file_next[5][27] ), .C(
        \reg_file_next[6][27] ), .D(\reg_file_next[7][27] ), .S0(n2231), .S1(
        n2215), .Y(n2893) );
  MXI4XL U2708 ( .A(\reg_file_next[20][27] ), .B(\reg_file_next[21][27] ), .C(
        \reg_file_next[22][27] ), .D(\reg_file_next[23][27] ), .S0(n2230), 
        .S1(n2214), .Y(n2889) );
  MXI4XL U2709 ( .A(\reg_file_next[4][28] ), .B(\reg_file_next[5][28] ), .C(
        \reg_file_next[6][28] ), .D(\reg_file_next[7][28] ), .S0(n2231), .S1(
        n2215), .Y(n2901) );
  MXI4XL U2710 ( .A(\reg_file_next[20][28] ), .B(\reg_file_next[21][28] ), .C(
        \reg_file_next[22][28] ), .D(\reg_file_next[23][28] ), .S0(n2231), 
        .S1(n2215), .Y(n2897) );
  MXI4XL U2711 ( .A(\reg_file_next[4][29] ), .B(\reg_file_next[5][29] ), .C(
        \reg_file_next[6][29] ), .D(\reg_file_next[7][29] ), .S0(n2232), .S1(
        n2215), .Y(n2909) );
  MXI4XL U2712 ( .A(\reg_file_next[20][29] ), .B(\reg_file_next[21][29] ), .C(
        \reg_file_next[22][29] ), .D(\reg_file_next[23][29] ), .S0(n2231), 
        .S1(n2215), .Y(n2905) );
  MXI4XL U2713 ( .A(\reg_file_next[4][30] ), .B(\reg_file_next[5][30] ), .C(
        \reg_file_next[6][30] ), .D(\reg_file_next[7][30] ), .S0(n2232), .S1(
        n2216), .Y(n2917) );
  MXI4XL U2714 ( .A(\reg_file_next[20][30] ), .B(\reg_file_next[21][30] ), .C(
        \reg_file_next[22][30] ), .D(\reg_file_next[23][30] ), .S0(n2232), 
        .S1(n2216), .Y(n2913) );
  MXI4XL U2715 ( .A(\reg_file_next[4][31] ), .B(\reg_file_next[5][31] ), .C(
        \reg_file_next[6][31] ), .D(\reg_file_next[7][31] ), .S0(n2233), .S1(
        n2216), .Y(n2925) );
  MXI4XL U2716 ( .A(\reg_file_next[20][31] ), .B(\reg_file_next[21][31] ), .C(
        \reg_file_next[22][31] ), .D(\reg_file_next[23][31] ), .S0(n2233), 
        .S1(n2216), .Y(n2921) );
  MXI4XL U2717 ( .A(\reg_file_next[4][0] ), .B(\reg_file_next[5][0] ), .C(
        \reg_file_next[6][0] ), .D(\reg_file_next[7][0] ), .S0(n2262), .S1(
        n2252), .Y(n2357) );
  MXI4XL U2718 ( .A(\reg_file_next[20][0] ), .B(\reg_file_next[21][0] ), .C(
        \reg_file_next[22][0] ), .D(\reg_file_next[23][0] ), .S0(n2262), .S1(
        n2252), .Y(n2353) );
  MXI4XL U2719 ( .A(\reg_file_next[4][1] ), .B(\reg_file_next[5][1] ), .C(
        \reg_file_next[6][1] ), .D(\reg_file_next[7][1] ), .S0(n2263), .S1(
        n2247), .Y(n2365) );
  MXI4XL U2720 ( .A(\reg_file_next[20][1] ), .B(\reg_file_next[21][1] ), .C(
        \reg_file_next[22][1] ), .D(\reg_file_next[23][1] ), .S0(n2263), .S1(
        n2252), .Y(n2361) );
  MXI4XL U2721 ( .A(\reg_file_next[4][2] ), .B(\reg_file_next[5][2] ), .C(
        \reg_file_next[6][2] ), .D(\reg_file_next[7][2] ), .S0(n2263), .S1(
        n2247), .Y(n2373) );
  MXI4XL U2722 ( .A(\reg_file_next[20][2] ), .B(\reg_file_next[21][2] ), .C(
        \reg_file_next[22][2] ), .D(\reg_file_next[23][2] ), .S0(n2263), .S1(
        n2247), .Y(n2369) );
  MXI4XL U2723 ( .A(\reg_file_next[4][3] ), .B(\reg_file_next[5][3] ), .C(
        \reg_file_next[6][3] ), .D(\reg_file_next[7][3] ), .S0(n2264), .S1(
        n2247), .Y(n2381) );
  MXI4XL U2724 ( .A(\reg_file_next[20][3] ), .B(\reg_file_next[21][3] ), .C(
        \reg_file_next[22][3] ), .D(\reg_file_next[23][3] ), .S0(n2264), .S1(
        n2247), .Y(n2377) );
  MXI4XL U2725 ( .A(\reg_file_next[4][4] ), .B(\reg_file_next[5][4] ), .C(
        \reg_file_next[6][4] ), .D(\reg_file_next[7][4] ), .S0(n2265), .S1(
        n2248), .Y(n2389) );
  MXI4XL U2726 ( .A(\reg_file_next[20][4] ), .B(\reg_file_next[21][4] ), .C(
        \reg_file_next[22][4] ), .D(\reg_file_next[23][4] ), .S0(n2264), .S1(
        n2248), .Y(n2385) );
  MXI4XL U2727 ( .A(\reg_file_next[4][5] ), .B(\reg_file_next[5][5] ), .C(
        \reg_file_next[6][5] ), .D(\reg_file_next[7][5] ), .S0(n2265), .S1(
        n2248), .Y(n2397) );
  MXI4XL U2728 ( .A(\reg_file_next[20][5] ), .B(\reg_file_next[21][5] ), .C(
        \reg_file_next[22][5] ), .D(\reg_file_next[23][5] ), .S0(n2265), .S1(
        n2248), .Y(n2393) );
  MXI4XL U2729 ( .A(\reg_file_next[4][6] ), .B(\reg_file_next[5][6] ), .C(
        \reg_file_next[6][6] ), .D(\reg_file_next[7][6] ), .S0(n2266), .S1(
        n2248), .Y(n2405) );
  MXI4XL U2730 ( .A(\reg_file_next[20][6] ), .B(\reg_file_next[21][6] ), .C(
        \reg_file_next[22][6] ), .D(\reg_file_next[23][6] ), .S0(n2265), .S1(
        n2248), .Y(n2401) );
  MXI4XL U2731 ( .A(\reg_file_next[4][7] ), .B(\reg_file_next[5][7] ), .C(
        \reg_file_next[6][7] ), .D(\reg_file_next[7][7] ), .S0(n2266), .S1(
        n2249), .Y(n2413) );
  MXI4XL U2732 ( .A(\reg_file_next[20][7] ), .B(\reg_file_next[21][7] ), .C(
        \reg_file_next[22][7] ), .D(\reg_file_next[23][7] ), .S0(n2266), .S1(
        n2249), .Y(n2409) );
  MXI4XL U2733 ( .A(\reg_file_next[4][8] ), .B(\reg_file_next[5][8] ), .C(
        \reg_file_next[6][8] ), .D(\reg_file_next[7][8] ), .S0(n2267), .S1(
        n2249), .Y(n2421) );
  MXI4XL U2734 ( .A(\reg_file_next[20][8] ), .B(\reg_file_next[21][8] ), .C(
        \reg_file_next[22][8] ), .D(\reg_file_next[23][8] ), .S0(n2267), .S1(
        n2249), .Y(n2417) );
  MXI4XL U2735 ( .A(\reg_file_next[4][9] ), .B(\reg_file_next[5][9] ), .C(
        \reg_file_next[6][9] ), .D(\reg_file_next[7][9] ), .S0(n2268), .S1(
        n2250), .Y(n2429) );
  MXI4XL U2736 ( .A(\reg_file_next[20][9] ), .B(\reg_file_next[21][9] ), .C(
        \reg_file_next[22][9] ), .D(\reg_file_next[23][9] ), .S0(n2267), .S1(
        n2249), .Y(n2425) );
  MXI4XL U2737 ( .A(\reg_file_next[4][10] ), .B(\reg_file_next[5][10] ), .C(
        \reg_file_next[6][10] ), .D(\reg_file_next[7][10] ), .S0(n2268), .S1(
        n2250), .Y(n2437) );
  MXI4XL U2738 ( .A(\reg_file_next[20][10] ), .B(\reg_file_next[21][10] ), .C(
        \reg_file_next[22][10] ), .D(\reg_file_next[23][10] ), .S0(n2268), 
        .S1(n2250), .Y(n2433) );
  MXI4XL U2739 ( .A(\reg_file_next[4][11] ), .B(\reg_file_next[5][11] ), .C(
        \reg_file_next[6][11] ), .D(\reg_file_next[7][11] ), .S0(n2269), .S1(
        n2250), .Y(n2445) );
  MXI4XL U2740 ( .A(\reg_file_next[20][11] ), .B(\reg_file_next[21][11] ), .C(
        \reg_file_next[22][11] ), .D(\reg_file_next[23][11] ), .S0(n2268), 
        .S1(n2250), .Y(n2441) );
  MXI4XL U2741 ( .A(\reg_file_next[4][12] ), .B(\reg_file_next[5][12] ), .C(
        \reg_file_next[6][12] ), .D(\reg_file_next[7][12] ), .S0(n2269), .S1(
        n2251), .Y(n2453) );
  MXI4XL U2742 ( .A(\reg_file_next[20][12] ), .B(\reg_file_next[21][12] ), .C(
        \reg_file_next[22][12] ), .D(\reg_file_next[23][12] ), .S0(n2269), 
        .S1(n2251), .Y(n2449) );
  MXI4XL U2743 ( .A(\reg_file_next[4][13] ), .B(\reg_file_next[5][13] ), .C(
        \reg_file_next[6][13] ), .D(\reg_file_next[7][13] ), .S0(n2270), .S1(
        n2251), .Y(n2461) );
  MXI4XL U2744 ( .A(\reg_file_next[20][13] ), .B(\reg_file_next[21][13] ), .C(
        \reg_file_next[22][13] ), .D(\reg_file_next[23][13] ), .S0(n2270), 
        .S1(n2251), .Y(n2457) );
  MXI4XL U2745 ( .A(\reg_file_next[4][14] ), .B(\reg_file_next[5][14] ), .C(
        \reg_file_next[6][14] ), .D(\reg_file_next[7][14] ), .S0(n2270), .S1(
        n2252), .Y(n2469) );
  MXI4XL U2746 ( .A(\reg_file_next[20][14] ), .B(\reg_file_next[21][14] ), .C(
        \reg_file_next[22][14] ), .D(\reg_file_next[23][14] ), .S0(n2270), 
        .S1(n2251), .Y(n2465) );
  MXI4XL U2747 ( .A(\reg_file_next[4][15] ), .B(\reg_file_next[5][15] ), .C(
        \reg_file_next[6][15] ), .D(\reg_file_next[7][15] ), .S0(n2259), .S1(
        n2252), .Y(n2477) );
  MXI4XL U2748 ( .A(\reg_file_next[20][15] ), .B(\reg_file_next[21][15] ), .C(
        \reg_file_next[22][15] ), .D(\reg_file_next[23][15] ), .S0(n2265), 
        .S1(n2252), .Y(n2473) );
  MXI4XL U2749 ( .A(\reg_file_next[4][16] ), .B(\reg_file_next[5][16] ), .C(
        \reg_file_next[6][16] ), .D(\reg_file_next[7][16] ), .S0(n2253), .S1(
        n2242), .Y(n2485) );
  MXI4XL U2750 ( .A(\reg_file_next[20][16] ), .B(\reg_file_next[21][16] ), .C(
        \reg_file_next[22][16] ), .D(\reg_file_next[23][16] ), .S0(n2253), 
        .S1(n2242), .Y(n2481) );
  MXI4XL U2751 ( .A(\reg_file_next[4][17] ), .B(\reg_file_next[5][17] ), .C(
        \reg_file_next[6][17] ), .D(\reg_file_next[7][17] ), .S0(n2254), .S1(
        n2243), .Y(n2493) );
  MXI4XL U2752 ( .A(\reg_file_next[20][17] ), .B(\reg_file_next[21][17] ), .C(
        \reg_file_next[22][17] ), .D(\reg_file_next[23][17] ), .S0(n2254), 
        .S1(n2242), .Y(n2489) );
  MXI4XL U2753 ( .A(\reg_file_next[4][18] ), .B(\reg_file_next[5][18] ), .C(
        \reg_file_next[6][18] ), .D(\reg_file_next[7][18] ), .S0(n2254), .S1(
        n2243), .Y(n2501) );
  MXI4XL U2754 ( .A(\reg_file_next[20][18] ), .B(\reg_file_next[21][18] ), .C(
        \reg_file_next[22][18] ), .D(\reg_file_next[23][18] ), .S0(n2254), 
        .S1(n2243), .Y(n2497) );
  MXI4XL U2755 ( .A(\reg_file_next[4][19] ), .B(\reg_file_next[5][19] ), .C(
        \reg_file_next[6][19] ), .D(\reg_file_next[7][19] ), .S0(n2255), .S1(
        n2243), .Y(n2509) );
  MXI4XL U2756 ( .A(\reg_file_next[20][19] ), .B(\reg_file_next[21][19] ), .C(
        \reg_file_next[22][19] ), .D(\reg_file_next[23][19] ), .S0(n2255), 
        .S1(n2243), .Y(n2505) );
  MXI4XL U2757 ( .A(\reg_file_next[4][20] ), .B(\reg_file_next[5][20] ), .C(
        \reg_file_next[6][20] ), .D(\reg_file_next[7][20] ), .S0(n2256), .S1(
        n2252), .Y(n2517) );
  MXI4XL U2758 ( .A(\reg_file_next[20][20] ), .B(\reg_file_next[21][20] ), .C(
        \reg_file_next[22][20] ), .D(\reg_file_next[23][20] ), .S0(n2255), 
        .S1(n2243), .Y(n2513) );
  MXI4XL U2759 ( .A(\reg_file_next[4][21] ), .B(\reg_file_next[5][21] ), .C(
        \reg_file_next[6][21] ), .D(\reg_file_next[7][21] ), .S0(n2256), .S1(
        n2243), .Y(n2525) );
  MXI4XL U2760 ( .A(\reg_file_next[20][21] ), .B(\reg_file_next[21][21] ), .C(
        \reg_file_next[22][21] ), .D(\reg_file_next[23][21] ), .S0(n2256), 
        .S1(n2247), .Y(n2521) );
  MXI4XL U2761 ( .A(\reg_file_next[4][22] ), .B(\reg_file_next[5][22] ), .C(
        \reg_file_next[6][22] ), .D(\reg_file_next[7][22] ), .S0(n2257), .S1(
        n2245), .Y(n2533) );
  MXI4XL U2762 ( .A(\reg_file_next[20][22] ), .B(\reg_file_next[21][22] ), .C(
        \reg_file_next[22][22] ), .D(\reg_file_next[23][22] ), .S0(n2256), 
        .S1(n2249), .Y(n2529) );
  MXI4XL U2763 ( .A(\reg_file_next[4][23] ), .B(\reg_file_next[5][23] ), .C(
        \reg_file_next[6][23] ), .D(\reg_file_next[7][23] ), .S0(n2257), .S1(
        n2244), .Y(n2541) );
  MXI4XL U2764 ( .A(\reg_file_next[20][23] ), .B(\reg_file_next[21][23] ), .C(
        \reg_file_next[22][23] ), .D(\reg_file_next[23][23] ), .S0(n2257), 
        .S1(n2244), .Y(n2537) );
  MXI4XL U2765 ( .A(\reg_file_next[4][24] ), .B(\reg_file_next[5][24] ), .C(
        \reg_file_next[6][24] ), .D(\reg_file_next[7][24] ), .S0(n2258), .S1(
        n2244), .Y(n2549) );
  MXI4XL U2766 ( .A(\reg_file_next[20][24] ), .B(\reg_file_next[21][24] ), .C(
        \reg_file_next[22][24] ), .D(\reg_file_next[23][24] ), .S0(n2258), 
        .S1(n2244), .Y(n2545) );
  MXI4XL U2767 ( .A(\reg_file_next[4][25] ), .B(\reg_file_next[5][25] ), .C(
        \reg_file_next[6][25] ), .D(\reg_file_next[7][25] ), .S0(n2258), .S1(
        n2245), .Y(n2557) );
  MXI4XL U2768 ( .A(\reg_file_next[20][25] ), .B(\reg_file_next[21][25] ), .C(
        \reg_file_next[22][25] ), .D(\reg_file_next[23][25] ), .S0(n2258), 
        .S1(n2244), .Y(n2553) );
  MXI4XL U2769 ( .A(\reg_file_next[4][26] ), .B(\reg_file_next[5][26] ), .C(
        \reg_file_next[6][26] ), .D(\reg_file_next[7][26] ), .S0(n2259), .S1(
        n2245), .Y(n2565) );
  MXI4XL U2770 ( .A(\reg_file_next[20][26] ), .B(\reg_file_next[21][26] ), .C(
        \reg_file_next[22][26] ), .D(\reg_file_next[23][26] ), .S0(n2259), 
        .S1(n2245), .Y(n2561) );
  MXI4XL U2771 ( .A(\reg_file_next[4][27] ), .B(\reg_file_next[5][27] ), .C(
        \reg_file_next[6][27] ), .D(\reg_file_next[7][27] ), .S0(n2260), .S1(
        n2245), .Y(n2573) );
  MXI4XL U2772 ( .A(\reg_file_next[20][27] ), .B(\reg_file_next[21][27] ), .C(
        \reg_file_next[22][27] ), .D(\reg_file_next[23][27] ), .S0(n2259), 
        .S1(n2245), .Y(n2569) );
  MXI4XL U2773 ( .A(\reg_file_next[4][28] ), .B(\reg_file_next[5][28] ), .C(
        \reg_file_next[6][28] ), .D(\reg_file_next[7][28] ), .S0(n2260), .S1(
        n2246), .Y(n2581) );
  MXI4XL U2774 ( .A(\reg_file_next[20][28] ), .B(\reg_file_next[21][28] ), .C(
        \reg_file_next[22][28] ), .D(\reg_file_next[23][28] ), .S0(n2260), 
        .S1(n2246), .Y(n2577) );
  MXI4XL U2775 ( .A(\reg_file_next[4][29] ), .B(\reg_file_next[5][29] ), .C(
        \reg_file_next[6][29] ), .D(\reg_file_next[7][29] ), .S0(n2261), .S1(
        n2246), .Y(n2589) );
  MXI4XL U2776 ( .A(\reg_file_next[20][29] ), .B(\reg_file_next[21][29] ), .C(
        \reg_file_next[22][29] ), .D(\reg_file_next[23][29] ), .S0(n2260), 
        .S1(n2246), .Y(n2585) );
  MXI4XL U2777 ( .A(\reg_file_next[4][30] ), .B(\reg_file_next[5][30] ), .C(
        \reg_file_next[6][30] ), .D(\reg_file_next[7][30] ), .S0(n2261), .S1(
        n2246), .Y(n2597) );
  MXI4XL U2778 ( .A(\reg_file_next[20][30] ), .B(\reg_file_next[21][30] ), .C(
        \reg_file_next[22][30] ), .D(\reg_file_next[23][30] ), .S0(n2261), 
        .S1(n2246), .Y(n2593) );
  MXI4XL U2779 ( .A(\reg_file_next[4][31] ), .B(\reg_file_next[5][31] ), .C(
        \reg_file_next[6][31] ), .D(\reg_file_next[7][31] ), .S0(n2262), .S1(
        n2242), .Y(n2605) );
  MXI4XL U2780 ( .A(\reg_file_next[20][31] ), .B(\reg_file_next[21][31] ), .C(
        \reg_file_next[22][31] ), .D(\reg_file_next[23][31] ), .S0(n2262), 
        .S1(n2245), .Y(n2601) );
  MXI4XL U2781 ( .A(\reg_file_next[0][0] ), .B(\reg_file_next[1][0] ), .C(
        \reg_file_next[2][0] ), .D(\reg_file_next[3][0] ), .S0(n2233), .S1(
        n2217), .Y(n2678) );
  MXI4XL U2782 ( .A(\reg_file_next[16][0] ), .B(\reg_file_next[17][0] ), .C(
        \reg_file_next[18][0] ), .D(\reg_file_next[19][0] ), .S0(n2233), .S1(
        n2216), .Y(n2674) );
  MXI4XL U2783 ( .A(\reg_file_next[0][1] ), .B(\reg_file_next[1][1] ), .C(
        \reg_file_next[2][1] ), .D(\reg_file_next[3][1] ), .S0(n2234), .S1(
        n2217), .Y(n2686) );
  MXI4XL U2784 ( .A(\reg_file_next[16][1] ), .B(\reg_file_next[17][1] ), .C(
        \reg_file_next[18][1] ), .D(\reg_file_next[19][1] ), .S0(n2234), .S1(
        n2217), .Y(n2682) );
  MXI4XL U2785 ( .A(\reg_file_next[0][2] ), .B(\reg_file_next[1][2] ), .C(
        \reg_file_next[2][2] ), .D(\reg_file_next[3][2] ), .S0(n2235), .S1(
        n2217), .Y(n2694) );
  MXI4XL U2786 ( .A(\reg_file_next[16][2] ), .B(\reg_file_next[17][2] ), .C(
        \reg_file_next[18][2] ), .D(\reg_file_next[19][2] ), .S0(n2234), .S1(
        n2217), .Y(n2690) );
  MXI4XL U2787 ( .A(\reg_file_next[0][3] ), .B(\reg_file_next[1][3] ), .C(
        \reg_file_next[2][3] ), .D(\reg_file_next[3][3] ), .S0(n2235), .S1(
        n2218), .Y(n2702) );
  MXI4XL U2788 ( .A(\reg_file_next[16][3] ), .B(\reg_file_next[17][3] ), .C(
        \reg_file_next[18][3] ), .D(\reg_file_next[19][3] ), .S0(n2235), .S1(
        n2218), .Y(n2698) );
  MXI4XL U2789 ( .A(\reg_file_next[0][4] ), .B(\reg_file_next[1][4] ), .C(
        \reg_file_next[2][4] ), .D(\reg_file_next[3][4] ), .S0(n2236), .S1(
        n2218), .Y(n2710) );
  MXI4XL U2790 ( .A(\reg_file_next[16][4] ), .B(\reg_file_next[17][4] ), .C(
        \reg_file_next[18][4] ), .D(\reg_file_next[19][4] ), .S0(n2235), .S1(
        n2218), .Y(n2706) );
  MXI4XL U2791 ( .A(\reg_file_next[0][5] ), .B(\reg_file_next[1][5] ), .C(
        \reg_file_next[2][5] ), .D(\reg_file_next[3][5] ), .S0(n2236), .S1(
        n2219), .Y(n2718) );
  MXI4XL U2792 ( .A(\reg_file_next[16][5] ), .B(\reg_file_next[17][5] ), .C(
        \reg_file_next[18][5] ), .D(\reg_file_next[19][5] ), .S0(n2236), .S1(
        n2218), .Y(n2714) );
  MXI4XL U2793 ( .A(\reg_file_next[0][6] ), .B(\reg_file_next[1][6] ), .C(
        \reg_file_next[2][6] ), .D(\reg_file_next[3][6] ), .S0(n2237), .S1(
        n2219), .Y(n2726) );
  MXI4XL U2794 ( .A(\reg_file_next[16][6] ), .B(\reg_file_next[17][6] ), .C(
        \reg_file_next[18][6] ), .D(\reg_file_next[19][6] ), .S0(n2237), .S1(
        n2219), .Y(n2722) );
  MXI4XL U2795 ( .A(\reg_file_next[0][7] ), .B(\reg_file_next[1][7] ), .C(
        \reg_file_next[2][7] ), .D(\reg_file_next[3][7] ), .S0(n2237), .S1(
        n2219), .Y(n2734) );
  MXI4XL U2796 ( .A(\reg_file_next[16][7] ), .B(\reg_file_next[17][7] ), .C(
        \reg_file_next[18][7] ), .D(\reg_file_next[19][7] ), .S0(n2237), .S1(
        n2219), .Y(n2730) );
  MXI4XL U2797 ( .A(\reg_file_next[0][8] ), .B(\reg_file_next[1][8] ), .C(
        \reg_file_next[2][8] ), .D(\reg_file_next[3][8] ), .S0(n2238), .S1(
        n2220), .Y(n2742) );
  MXI4XL U2798 ( .A(\reg_file_next[16][8] ), .B(\reg_file_next[17][8] ), .C(
        \reg_file_next[18][8] ), .D(\reg_file_next[19][8] ), .S0(n2238), .S1(
        n2220), .Y(n2738) );
  MXI4XL U2799 ( .A(\reg_file_next[0][9] ), .B(\reg_file_next[1][9] ), .C(
        \reg_file_next[2][9] ), .D(\reg_file_next[3][9] ), .S0(n2239), .S1(
        n2220), .Y(n2750) );
  MXI4XL U2800 ( .A(\reg_file_next[16][9] ), .B(\reg_file_next[17][9] ), .C(
        \reg_file_next[18][9] ), .D(\reg_file_next[19][9] ), .S0(n2238), .S1(
        n2220), .Y(n2746) );
  MXI4XL U2801 ( .A(\reg_file_next[0][10] ), .B(\reg_file_next[1][10] ), .C(
        \reg_file_next[2][10] ), .D(\reg_file_next[3][10] ), .S0(n2239), .S1(
        n2221), .Y(n2758) );
  MXI4XL U2802 ( .A(\reg_file_next[16][10] ), .B(\reg_file_next[17][10] ), .C(
        \reg_file_next[18][10] ), .D(\reg_file_next[19][10] ), .S0(n2239), 
        .S1(n2220), .Y(n2754) );
  MXI4XL U2803 ( .A(\reg_file_next[0][11] ), .B(\reg_file_next[1][11] ), .C(
        \reg_file_next[2][11] ), .D(\reg_file_next[3][11] ), .S0(n2240), .S1(
        n2221), .Y(n2766) );
  MXI4XL U2804 ( .A(\reg_file_next[16][11] ), .B(\reg_file_next[17][11] ), .C(
        \reg_file_next[18][11] ), .D(\reg_file_next[19][11] ), .S0(n2239), 
        .S1(n2221), .Y(n2762) );
  MXI4XL U2805 ( .A(\reg_file_next[0][12] ), .B(\reg_file_next[1][12] ), .C(
        \reg_file_next[2][12] ), .D(\reg_file_next[3][12] ), .S0(n2240), .S1(
        n2221), .Y(n2774) );
  MXI4XL U2806 ( .A(\reg_file_next[16][12] ), .B(\reg_file_next[17][12] ), .C(
        \reg_file_next[18][12] ), .D(\reg_file_next[19][12] ), .S0(n2240), 
        .S1(n2221), .Y(n2770) );
  MXI4XL U2807 ( .A(\reg_file_next[0][13] ), .B(\reg_file_next[1][13] ), .C(
        \reg_file_next[2][13] ), .D(\reg_file_next[3][13] ), .S0(n2241), .S1(
        n2222), .Y(n2782) );
  MXI4XL U2808 ( .A(\reg_file_next[16][13] ), .B(\reg_file_next[17][13] ), .C(
        \reg_file_next[18][13] ), .D(\reg_file_next[19][13] ), .S0(n2241), 
        .S1(n2222), .Y(n2778) );
  MXI4XL U2809 ( .A(\reg_file_next[0][14] ), .B(\reg_file_next[1][14] ), .C(
        \reg_file_next[2][14] ), .D(\reg_file_next[3][14] ), .S0(n2241), .S1(
        n2222), .Y(n2790) );
  MXI4XL U2810 ( .A(\reg_file_next[16][14] ), .B(\reg_file_next[17][14] ), .C(
        \reg_file_next[18][14] ), .D(\reg_file_next[19][14] ), .S0(n2241), 
        .S1(n2222), .Y(n2786) );
  MXI4XL U2811 ( .A(\reg_file_next[0][15] ), .B(\reg_file_next[1][15] ), .C(
        \reg_file_next[2][15] ), .D(\reg_file_next[3][15] ), .S0(n2229), .S1(
        n2223), .Y(n2798) );
  MXI4XL U2812 ( .A(\reg_file_next[16][15] ), .B(\reg_file_next[17][15] ), .C(
        \reg_file_next[18][15] ), .D(\reg_file_next[19][15] ), .S0(n2236), 
        .S1(n2222), .Y(n2794) );
  MXI4XL U2813 ( .A(\reg_file_next[0][16] ), .B(\reg_file_next[1][16] ), .C(
        \reg_file_next[2][16] ), .D(\reg_file_next[3][16] ), .S0(n2224), .S1(
        n2210), .Y(n2806) );
  MXI4XL U2814 ( .A(\reg_file_next[16][16] ), .B(\reg_file_next[17][16] ), .C(
        \reg_file_next[18][16] ), .D(\reg_file_next[19][16] ), .S0(n2224), 
        .S1(n2210), .Y(n2802) );
  MXI4XL U2815 ( .A(\reg_file_next[0][17] ), .B(\reg_file_next[1][17] ), .C(
        \reg_file_next[2][17] ), .D(\reg_file_next[3][17] ), .S0(n2225), .S1(
        n2211), .Y(n2814) );
  MXI4XL U2816 ( .A(\reg_file_next[16][17] ), .B(\reg_file_next[17][17] ), .C(
        \reg_file_next[18][17] ), .D(\reg_file_next[19][17] ), .S0(n2225), 
        .S1(n2210), .Y(n2810) );
  MXI4XL U2817 ( .A(\reg_file_next[0][18] ), .B(\reg_file_next[1][18] ), .C(
        \reg_file_next[2][18] ), .D(\reg_file_next[3][18] ), .S0(n2225), .S1(
        n2211), .Y(n2822) );
  MXI4XL U2818 ( .A(\reg_file_next[16][18] ), .B(\reg_file_next[17][18] ), .C(
        \reg_file_next[18][18] ), .D(\reg_file_next[19][18] ), .S0(n2225), 
        .S1(n2211), .Y(n2818) );
  MXI4XL U2819 ( .A(\reg_file_next[0][19] ), .B(\reg_file_next[1][19] ), .C(
        \reg_file_next[2][19] ), .D(\reg_file_next[3][19] ), .S0(n2226), .S1(
        n2211), .Y(n2830) );
  MXI4XL U2820 ( .A(\reg_file_next[16][19] ), .B(\reg_file_next[17][19] ), .C(
        \reg_file_next[18][19] ), .D(\reg_file_next[19][19] ), .S0(n2226), 
        .S1(n2211), .Y(n2826) );
  MXI4XL U2821 ( .A(\reg_file_next[0][20] ), .B(\reg_file_next[1][20] ), .C(
        \reg_file_next[2][20] ), .D(\reg_file_next[3][20] ), .S0(n2227), .S1(
        n2212), .Y(n2838) );
  MXI4XL U2822 ( .A(\reg_file_next[16][20] ), .B(\reg_file_next[17][20] ), .C(
        \reg_file_next[18][20] ), .D(\reg_file_next[19][20] ), .S0(n2226), 
        .S1(n2212), .Y(n2834) );
  MXI4XL U2823 ( .A(\reg_file_next[0][21] ), .B(\reg_file_next[1][21] ), .C(
        \reg_file_next[2][21] ), .D(\reg_file_next[3][21] ), .S0(n2227), .S1(
        n2212), .Y(n2846) );
  MXI4XL U2824 ( .A(\reg_file_next[16][21] ), .B(\reg_file_next[17][21] ), .C(
        \reg_file_next[18][21] ), .D(\reg_file_next[19][21] ), .S0(n2227), 
        .S1(n2212), .Y(n2842) );
  MXI4XL U2825 ( .A(\reg_file_next[0][22] ), .B(\reg_file_next[1][22] ), .C(
        \reg_file_next[2][22] ), .D(\reg_file_next[3][22] ), .S0(n2228), .S1(
        n2213), .Y(n2854) );
  MXI4XL U2826 ( .A(\reg_file_next[16][22] ), .B(\reg_file_next[17][22] ), .C(
        \reg_file_next[18][22] ), .D(\reg_file_next[19][22] ), .S0(n2227), 
        .S1(n2212), .Y(n2850) );
  MXI4XL U2827 ( .A(\reg_file_next[0][23] ), .B(\reg_file_next[1][23] ), .C(
        \reg_file_next[2][23] ), .D(\reg_file_next[3][23] ), .S0(n2228), .S1(
        n2213), .Y(n2862) );
  MXI4XL U2828 ( .A(\reg_file_next[16][23] ), .B(\reg_file_next[17][23] ), .C(
        \reg_file_next[18][23] ), .D(\reg_file_next[19][23] ), .S0(n2228), 
        .S1(n2213), .Y(n2858) );
  MXI4XL U2829 ( .A(\reg_file_next[0][24] ), .B(\reg_file_next[1][24] ), .C(
        \reg_file_next[2][24] ), .D(\reg_file_next[3][24] ), .S0(n2229), .S1(
        n2213), .Y(n2870) );
  MXI4XL U2830 ( .A(\reg_file_next[16][24] ), .B(\reg_file_next[17][24] ), .C(
        \reg_file_next[18][24] ), .D(\reg_file_next[19][24] ), .S0(n2229), 
        .S1(n2213), .Y(n2866) );
  MXI4XL U2831 ( .A(\reg_file_next[0][25] ), .B(\reg_file_next[1][25] ), .C(
        \reg_file_next[2][25] ), .D(\reg_file_next[3][25] ), .S0(n2229), .S1(
        n2214), .Y(n2878) );
  MXI4XL U2832 ( .A(\reg_file_next[16][25] ), .B(\reg_file_next[17][25] ), .C(
        \reg_file_next[18][25] ), .D(\reg_file_next[19][25] ), .S0(n2229), 
        .S1(n2214), .Y(n2874) );
  MXI4XL U2833 ( .A(\reg_file_next[0][26] ), .B(\reg_file_next[1][26] ), .C(
        \reg_file_next[2][26] ), .D(\reg_file_next[3][26] ), .S0(n2230), .S1(
        n2214), .Y(n2886) );
  MXI4XL U2834 ( .A(\reg_file_next[16][26] ), .B(\reg_file_next[17][26] ), .C(
        \reg_file_next[18][26] ), .D(\reg_file_next[19][26] ), .S0(n2230), 
        .S1(n2214), .Y(n2882) );
  MXI4XL U2835 ( .A(\reg_file_next[0][27] ), .B(\reg_file_next[1][27] ), .C(
        \reg_file_next[2][27] ), .D(\reg_file_next[3][27] ), .S0(n2231), .S1(
        n2215), .Y(n2894) );
  MXI4XL U2836 ( .A(\reg_file_next[16][27] ), .B(\reg_file_next[17][27] ), .C(
        \reg_file_next[18][27] ), .D(\reg_file_next[19][27] ), .S0(n2230), 
        .S1(n2214), .Y(n2890) );
  MXI4XL U2837 ( .A(\reg_file_next[0][28] ), .B(\reg_file_next[1][28] ), .C(
        \reg_file_next[2][28] ), .D(\reg_file_next[3][28] ), .S0(n2231), .S1(
        n2215), .Y(n2902) );
  MXI4XL U2838 ( .A(\reg_file_next[16][28] ), .B(\reg_file_next[17][28] ), .C(
        \reg_file_next[18][28] ), .D(\reg_file_next[19][28] ), .S0(n2231), 
        .S1(n2215), .Y(n2898) );
  MXI4XL U2839 ( .A(\reg_file_next[0][29] ), .B(\reg_file_next[1][29] ), .C(
        \reg_file_next[2][29] ), .D(\reg_file_next[3][29] ), .S0(n2232), .S1(
        n2215), .Y(n2910) );
  MXI4XL U2840 ( .A(\reg_file_next[16][29] ), .B(\reg_file_next[17][29] ), .C(
        \reg_file_next[18][29] ), .D(\reg_file_next[19][29] ), .S0(n2231), 
        .S1(n2215), .Y(n2906) );
  MXI4XL U2841 ( .A(\reg_file_next[0][30] ), .B(\reg_file_next[1][30] ), .C(
        \reg_file_next[2][30] ), .D(\reg_file_next[3][30] ), .S0(n2232), .S1(
        n2216), .Y(n2918) );
  MXI4XL U2842 ( .A(\reg_file_next[16][30] ), .B(\reg_file_next[17][30] ), .C(
        \reg_file_next[18][30] ), .D(\reg_file_next[19][30] ), .S0(n2232), 
        .S1(n2216), .Y(n2914) );
  MXI4XL U2843 ( .A(\reg_file_next[0][31] ), .B(\reg_file_next[1][31] ), .C(
        \reg_file_next[2][31] ), .D(\reg_file_next[3][31] ), .S0(n2233), .S1(
        n2216), .Y(n2926) );
  MXI4XL U2844 ( .A(\reg_file_next[16][31] ), .B(\reg_file_next[17][31] ), .C(
        \reg_file_next[18][31] ), .D(\reg_file_next[19][31] ), .S0(n2233), 
        .S1(n2216), .Y(n2922) );
  MXI4XL U2845 ( .A(\reg_file_next[0][0] ), .B(\reg_file_next[1][0] ), .C(
        \reg_file_next[2][0] ), .D(\reg_file_next[3][0] ), .S0(n2262), .S1(
        n2249), .Y(n2358) );
  MXI4XL U2846 ( .A(\reg_file_next[16][0] ), .B(\reg_file_next[17][0] ), .C(
        \reg_file_next[18][0] ), .D(\reg_file_next[19][0] ), .S0(n2262), .S1(
        n2246), .Y(n2354) );
  MXI4XL U2847 ( .A(\reg_file_next[0][1] ), .B(\reg_file_next[1][1] ), .C(
        \reg_file_next[2][1] ), .D(\reg_file_next[3][1] ), .S0(n2263), .S1(
        n2247), .Y(n2366) );
  MXI4XL U2848 ( .A(\reg_file_next[16][1] ), .B(\reg_file_next[17][1] ), .C(
        \reg_file_next[18][1] ), .D(\reg_file_next[19][1] ), .S0(n2263), .S1(
        n2244), .Y(n2362) );
  MXI4XL U2849 ( .A(\reg_file_next[0][2] ), .B(\reg_file_next[1][2] ), .C(
        \reg_file_next[2][2] ), .D(\reg_file_next[3][2] ), .S0(n2264), .S1(
        n2247), .Y(n2374) );
  MXI4XL U2850 ( .A(\reg_file_next[16][2] ), .B(\reg_file_next[17][2] ), .C(
        \reg_file_next[18][2] ), .D(\reg_file_next[19][2] ), .S0(n2263), .S1(
        n2247), .Y(n2370) );
  MXI4XL U2851 ( .A(\reg_file_next[0][3] ), .B(\reg_file_next[1][3] ), .C(
        \reg_file_next[2][3] ), .D(\reg_file_next[3][3] ), .S0(n2264), .S1(
        n2247), .Y(n2382) );
  MXI4XL U2852 ( .A(\reg_file_next[16][3] ), .B(\reg_file_next[17][3] ), .C(
        \reg_file_next[18][3] ), .D(\reg_file_next[19][3] ), .S0(n2264), .S1(
        n2247), .Y(n2378) );
  MXI4XL U2853 ( .A(\reg_file_next[0][4] ), .B(\reg_file_next[1][4] ), .C(
        \reg_file_next[2][4] ), .D(\reg_file_next[3][4] ), .S0(n2265), .S1(
        n2248), .Y(n2390) );
  MXI4XL U2854 ( .A(\reg_file_next[16][4] ), .B(\reg_file_next[17][4] ), .C(
        \reg_file_next[18][4] ), .D(\reg_file_next[19][4] ), .S0(n2264), .S1(
        n2248), .Y(n2386) );
  MXI4XL U2855 ( .A(\reg_file_next[0][5] ), .B(\reg_file_next[1][5] ), .C(
        \reg_file_next[2][5] ), .D(\reg_file_next[3][5] ), .S0(n2265), .S1(
        n2248), .Y(n2398) );
  MXI4XL U2856 ( .A(\reg_file_next[16][5] ), .B(\reg_file_next[17][5] ), .C(
        \reg_file_next[18][5] ), .D(\reg_file_next[19][5] ), .S0(n2265), .S1(
        n2248), .Y(n2394) );
  MXI4XL U2857 ( .A(\reg_file_next[0][6] ), .B(\reg_file_next[1][6] ), .C(
        \reg_file_next[2][6] ), .D(\reg_file_next[3][6] ), .S0(n2266), .S1(
        n2249), .Y(n2406) );
  MXI4XL U2858 ( .A(\reg_file_next[16][6] ), .B(\reg_file_next[17][6] ), .C(
        \reg_file_next[18][6] ), .D(\reg_file_next[19][6] ), .S0(n2266), .S1(
        n2248), .Y(n2402) );
  MXI4XL U2859 ( .A(\reg_file_next[0][7] ), .B(\reg_file_next[1][7] ), .C(
        \reg_file_next[2][7] ), .D(\reg_file_next[3][7] ), .S0(n2266), .S1(
        n2249), .Y(n2414) );
  MXI4XL U2860 ( .A(\reg_file_next[16][7] ), .B(\reg_file_next[17][7] ), .C(
        \reg_file_next[18][7] ), .D(\reg_file_next[19][7] ), .S0(n2266), .S1(
        n2249), .Y(n2410) );
  MXI4XL U2861 ( .A(\reg_file_next[0][8] ), .B(\reg_file_next[1][8] ), .C(
        \reg_file_next[2][8] ), .D(\reg_file_next[3][8] ), .S0(n2267), .S1(
        n2249), .Y(n2422) );
  MXI4XL U2862 ( .A(\reg_file_next[16][8] ), .B(\reg_file_next[17][8] ), .C(
        \reg_file_next[18][8] ), .D(\reg_file_next[19][8] ), .S0(n2267), .S1(
        n2249), .Y(n2418) );
  MXI4XL U2863 ( .A(\reg_file_next[0][9] ), .B(\reg_file_next[1][9] ), .C(
        \reg_file_next[2][9] ), .D(\reg_file_next[3][9] ), .S0(n2268), .S1(
        n2250), .Y(n2430) );
  MXI4XL U2864 ( .A(\reg_file_next[16][9] ), .B(\reg_file_next[17][9] ), .C(
        \reg_file_next[18][9] ), .D(\reg_file_next[19][9] ), .S0(n2267), .S1(
        n2250), .Y(n2426) );
  MXI4XL U2865 ( .A(\reg_file_next[0][10] ), .B(\reg_file_next[1][10] ), .C(
        \reg_file_next[2][10] ), .D(\reg_file_next[3][10] ), .S0(n2268), .S1(
        n2250), .Y(n2438) );
  MXI4XL U2866 ( .A(\reg_file_next[16][10] ), .B(\reg_file_next[17][10] ), .C(
        \reg_file_next[18][10] ), .D(\reg_file_next[19][10] ), .S0(n2268), 
        .S1(n2250), .Y(n2434) );
  MXI4XL U2867 ( .A(\reg_file_next[0][11] ), .B(\reg_file_next[1][11] ), .C(
        \reg_file_next[2][11] ), .D(\reg_file_next[3][11] ), .S0(n2269), .S1(
        n2250), .Y(n2446) );
  MXI4XL U2868 ( .A(\reg_file_next[16][11] ), .B(\reg_file_next[17][11] ), .C(
        \reg_file_next[18][11] ), .D(\reg_file_next[19][11] ), .S0(n2268), 
        .S1(n2250), .Y(n2442) );
  MXI4XL U2869 ( .A(\reg_file_next[0][12] ), .B(\reg_file_next[1][12] ), .C(
        \reg_file_next[2][12] ), .D(\reg_file_next[3][12] ), .S0(n2269), .S1(
        n2251), .Y(n2454) );
  MXI4XL U2870 ( .A(\reg_file_next[16][12] ), .B(\reg_file_next[17][12] ), .C(
        \reg_file_next[18][12] ), .D(\reg_file_next[19][12] ), .S0(n2269), 
        .S1(n2251), .Y(n2450) );
  MXI4XL U2871 ( .A(\reg_file_next[0][13] ), .B(\reg_file_next[1][13] ), .C(
        \reg_file_next[2][13] ), .D(\reg_file_next[3][13] ), .S0(n2270), .S1(
        n2251), .Y(n2462) );
  MXI4XL U2872 ( .A(\reg_file_next[16][13] ), .B(\reg_file_next[17][13] ), .C(
        \reg_file_next[18][13] ), .D(\reg_file_next[19][13] ), .S0(n2270), 
        .S1(n2251), .Y(n2458) );
  MXI4XL U2873 ( .A(\reg_file_next[0][14] ), .B(\reg_file_next[1][14] ), .C(
        \reg_file_next[2][14] ), .D(\reg_file_next[3][14] ), .S0(n2270), .S1(
        n2252), .Y(n2470) );
  MXI4XL U2874 ( .A(\reg_file_next[16][14] ), .B(\reg_file_next[17][14] ), .C(
        \reg_file_next[18][14] ), .D(\reg_file_next[19][14] ), .S0(n2270), 
        .S1(n2251), .Y(n2466) );
  MXI4XL U2875 ( .A(\reg_file_next[0][15] ), .B(\reg_file_next[1][15] ), .C(
        \reg_file_next[2][15] ), .D(\reg_file_next[3][15] ), .S0(n2263), .S1(
        n2252), .Y(n2478) );
  MXI4XL U2876 ( .A(\reg_file_next[16][15] ), .B(\reg_file_next[17][15] ), .C(
        \reg_file_next[18][15] ), .D(\reg_file_next[19][15] ), .S0(n2269), 
        .S1(n2252), .Y(n2474) );
  MXI4XL U2877 ( .A(\reg_file_next[0][16] ), .B(\reg_file_next[1][16] ), .C(
        \reg_file_next[2][16] ), .D(\reg_file_next[3][16] ), .S0(n2253), .S1(
        n2242), .Y(n2486) );
  MXI4XL U2878 ( .A(\reg_file_next[16][16] ), .B(\reg_file_next[17][16] ), .C(
        \reg_file_next[18][16] ), .D(\reg_file_next[19][16] ), .S0(n2253), 
        .S1(n2242), .Y(n2482) );
  MXI4XL U2879 ( .A(\reg_file_next[0][17] ), .B(\reg_file_next[1][17] ), .C(
        \reg_file_next[2][17] ), .D(\reg_file_next[3][17] ), .S0(n2254), .S1(
        n2243), .Y(n2494) );
  MXI4XL U2880 ( .A(\reg_file_next[16][17] ), .B(\reg_file_next[17][17] ), .C(
        \reg_file_next[18][17] ), .D(\reg_file_next[19][17] ), .S0(n2254), 
        .S1(n2242), .Y(n2490) );
  MXI4XL U2881 ( .A(\reg_file_next[0][18] ), .B(\reg_file_next[1][18] ), .C(
        \reg_file_next[2][18] ), .D(\reg_file_next[3][18] ), .S0(n2254), .S1(
        n2243), .Y(n2502) );
  MXI4XL U2882 ( .A(\reg_file_next[16][18] ), .B(\reg_file_next[17][18] ), .C(
        \reg_file_next[18][18] ), .D(\reg_file_next[19][18] ), .S0(n2254), 
        .S1(n2243), .Y(n2498) );
  MXI4XL U2883 ( .A(\reg_file_next[0][19] ), .B(\reg_file_next[1][19] ), .C(
        \reg_file_next[2][19] ), .D(\reg_file_next[3][19] ), .S0(n2255), .S1(
        n2243), .Y(n2510) );
  MXI4XL U2884 ( .A(\reg_file_next[16][19] ), .B(\reg_file_next[17][19] ), .C(
        \reg_file_next[18][19] ), .D(\reg_file_next[19][19] ), .S0(n2255), 
        .S1(n2243), .Y(n2506) );
  MXI4XL U2885 ( .A(\reg_file_next[0][20] ), .B(\reg_file_next[1][20] ), .C(
        \reg_file_next[2][20] ), .D(\reg_file_next[3][20] ), .S0(n2256), .S1(
        n2246), .Y(n2518) );
  MXI4XL U2886 ( .A(\reg_file_next[16][20] ), .B(\reg_file_next[17][20] ), .C(
        \reg_file_next[18][20] ), .D(\reg_file_next[19][20] ), .S0(n2255), 
        .S1(n2244), .Y(n2514) );
  MXI4XL U2887 ( .A(\reg_file_next[0][21] ), .B(\reg_file_next[1][21] ), .C(
        \reg_file_next[2][21] ), .D(\reg_file_next[3][21] ), .S0(n2256), .S1(
        n2250), .Y(n2526) );
  MXI4XL U2888 ( .A(\reg_file_next[16][21] ), .B(\reg_file_next[17][21] ), .C(
        \reg_file_next[18][21] ), .D(\reg_file_next[19][21] ), .S0(n2256), 
        .S1(n2248), .Y(n2522) );
  MXI4XL U2889 ( .A(\reg_file_next[0][22] ), .B(\reg_file_next[1][22] ), .C(
        \reg_file_next[2][22] ), .D(\reg_file_next[3][22] ), .S0(n2257), .S1(
        n2251), .Y(n2534) );
  MXI4XL U2890 ( .A(\reg_file_next[16][22] ), .B(\reg_file_next[17][22] ), .C(
        \reg_file_next[18][22] ), .D(\reg_file_next[19][22] ), .S0(n2256), 
        .S1(n2243), .Y(n2530) );
  MXI4XL U2891 ( .A(\reg_file_next[0][23] ), .B(\reg_file_next[1][23] ), .C(
        \reg_file_next[2][23] ), .D(\reg_file_next[3][23] ), .S0(n2257), .S1(
        n2244), .Y(n2542) );
  MXI4XL U2892 ( .A(\reg_file_next[16][23] ), .B(\reg_file_next[17][23] ), .C(
        \reg_file_next[18][23] ), .D(\reg_file_next[19][23] ), .S0(n2257), 
        .S1(n2244), .Y(n2538) );
  MXI4XL U2893 ( .A(\reg_file_next[0][24] ), .B(\reg_file_next[1][24] ), .C(
        \reg_file_next[2][24] ), .D(\reg_file_next[3][24] ), .S0(n2258), .S1(
        n2244), .Y(n2550) );
  MXI4XL U2894 ( .A(\reg_file_next[16][24] ), .B(\reg_file_next[17][24] ), .C(
        \reg_file_next[18][24] ), .D(\reg_file_next[19][24] ), .S0(n2258), 
        .S1(n2244), .Y(n2546) );
  MXI4XL U2895 ( .A(\reg_file_next[0][25] ), .B(\reg_file_next[1][25] ), .C(
        \reg_file_next[2][25] ), .D(\reg_file_next[3][25] ), .S0(n2258), .S1(
        n2245), .Y(n2558) );
  MXI4XL U2896 ( .A(\reg_file_next[16][25] ), .B(\reg_file_next[17][25] ), .C(
        \reg_file_next[18][25] ), .D(\reg_file_next[19][25] ), .S0(n2258), 
        .S1(n2244), .Y(n2554) );
  MXI4XL U2897 ( .A(\reg_file_next[0][26] ), .B(\reg_file_next[1][26] ), .C(
        \reg_file_next[2][26] ), .D(\reg_file_next[3][26] ), .S0(n2259), .S1(
        n2245), .Y(n2566) );
  MXI4XL U2898 ( .A(\reg_file_next[16][26] ), .B(\reg_file_next[17][26] ), .C(
        \reg_file_next[18][26] ), .D(\reg_file_next[19][26] ), .S0(n2259), 
        .S1(n2245), .Y(n2562) );
  MXI4XL U2899 ( .A(\reg_file_next[0][27] ), .B(\reg_file_next[1][27] ), .C(
        \reg_file_next[2][27] ), .D(\reg_file_next[3][27] ), .S0(n2260), .S1(
        n2245), .Y(n2574) );
  MXI4XL U2900 ( .A(\reg_file_next[16][27] ), .B(\reg_file_next[17][27] ), .C(
        \reg_file_next[18][27] ), .D(\reg_file_next[19][27] ), .S0(n2259), 
        .S1(n2245), .Y(n2570) );
  MXI4XL U2901 ( .A(\reg_file_next[0][28] ), .B(\reg_file_next[1][28] ), .C(
        \reg_file_next[2][28] ), .D(\reg_file_next[3][28] ), .S0(n2260), .S1(
        n2246), .Y(n2582) );
  MXI4XL U2902 ( .A(\reg_file_next[16][28] ), .B(\reg_file_next[17][28] ), .C(
        \reg_file_next[18][28] ), .D(\reg_file_next[19][28] ), .S0(n2260), 
        .S1(n2246), .Y(n2578) );
  MXI4XL U2903 ( .A(\reg_file_next[0][29] ), .B(\reg_file_next[1][29] ), .C(
        \reg_file_next[2][29] ), .D(\reg_file_next[3][29] ), .S0(n2261), .S1(
        n2246), .Y(n2590) );
  MXI4XL U2904 ( .A(\reg_file_next[16][29] ), .B(\reg_file_next[17][29] ), .C(
        \reg_file_next[18][29] ), .D(\reg_file_next[19][29] ), .S0(n2260), 
        .S1(n2246), .Y(n2586) );
  MXI4XL U2905 ( .A(\reg_file_next[0][30] ), .B(\reg_file_next[1][30] ), .C(
        \reg_file_next[2][30] ), .D(\reg_file_next[3][30] ), .S0(n2261), .S1(
        n2250), .Y(n2598) );
  MXI4XL U2906 ( .A(\reg_file_next[16][30] ), .B(\reg_file_next[17][30] ), .C(
        \reg_file_next[18][30] ), .D(\reg_file_next[19][30] ), .S0(n2261), 
        .S1(n2246), .Y(n2594) );
  MXI4XL U2907 ( .A(\reg_file_next[0][31] ), .B(\reg_file_next[1][31] ), .C(
        \reg_file_next[2][31] ), .D(\reg_file_next[3][31] ), .S0(n2262), .S1(
        n2248), .Y(n2606) );
  MXI4XL U2908 ( .A(\reg_file_next[16][31] ), .B(\reg_file_next[17][31] ), .C(
        \reg_file_next[18][31] ), .D(\reg_file_next[19][31] ), .S0(n2262), 
        .S1(n2251), .Y(n2602) );
  MXI4XL U2909 ( .A(\reg_file_next[12][0] ), .B(\reg_file_next[13][0] ), .C(
        \reg_file_next[14][0] ), .D(\reg_file_next[15][0] ), .S0(n2233), .S1(
        n2216), .Y(n2675) );
  MXI4XL U2910 ( .A(\reg_file_next[28][0] ), .B(\reg_file_next[29][0] ), .C(
        \reg_file_next[30][0] ), .D(\reg_file_next[31][0] ), .S0(n2224), .S1(
        n2210), .Y(n2671) );
  MXI4XL U2911 ( .A(\reg_file_next[12][1] ), .B(\reg_file_next[13][1] ), .C(
        \reg_file_next[14][1] ), .D(\reg_file_next[15][1] ), .S0(n2234), .S1(
        n2217), .Y(n2683) );
  MXI4XL U2912 ( .A(\reg_file_next[28][1] ), .B(\reg_file_next[29][1] ), .C(
        \reg_file_next[30][1] ), .D(\reg_file_next[31][1] ), .S0(n2233), .S1(
        n2217), .Y(n2679) );
  MXI4XL U2913 ( .A(\reg_file_next[12][2] ), .B(\reg_file_next[13][2] ), .C(
        \reg_file_next[14][2] ), .D(\reg_file_next[15][2] ), .S0(n2234), .S1(
        n2217), .Y(n2691) );
  MXI4XL U2914 ( .A(\reg_file_next[28][2] ), .B(\reg_file_next[29][2] ), .C(
        \reg_file_next[30][2] ), .D(\reg_file_next[31][2] ), .S0(n2234), .S1(
        n2217), .Y(n2687) );
  MXI4XL U2915 ( .A(\reg_file_next[12][3] ), .B(\reg_file_next[13][3] ), .C(
        \reg_file_next[14][3] ), .D(\reg_file_next[15][3] ), .S0(n2235), .S1(
        n2218), .Y(n2699) );
  MXI4XL U2916 ( .A(\reg_file_next[28][3] ), .B(\reg_file_next[29][3] ), .C(
        \reg_file_next[30][3] ), .D(\reg_file_next[31][3] ), .S0(n2235), .S1(
        n2217), .Y(n2695) );
  MXI4XL U2917 ( .A(\reg_file_next[12][4] ), .B(\reg_file_next[13][4] ), .C(
        \reg_file_next[14][4] ), .D(\reg_file_next[15][4] ), .S0(n2235), .S1(
        n2218), .Y(n2707) );
  MXI4XL U2918 ( .A(\reg_file_next[28][4] ), .B(\reg_file_next[29][4] ), .C(
        \reg_file_next[30][4] ), .D(\reg_file_next[31][4] ), .S0(n2235), .S1(
        n2218), .Y(n2703) );
  MXI4XL U2919 ( .A(\reg_file_next[12][5] ), .B(\reg_file_next[13][5] ), .C(
        \reg_file_next[14][5] ), .D(\reg_file_next[15][5] ), .S0(n2236), .S1(
        n2218), .Y(n2715) );
  MXI4XL U2920 ( .A(\reg_file_next[28][5] ), .B(\reg_file_next[29][5] ), .C(
        \reg_file_next[30][5] ), .D(\reg_file_next[31][5] ), .S0(n2236), .S1(
        n2218), .Y(n2711) );
  MXI4XL U2921 ( .A(\reg_file_next[12][6] ), .B(\reg_file_next[13][6] ), .C(
        \reg_file_next[14][6] ), .D(\reg_file_next[15][6] ), .S0(n2237), .S1(
        n2219), .Y(n2723) );
  MXI4XL U2922 ( .A(\reg_file_next[28][6] ), .B(\reg_file_next[29][6] ), .C(
        \reg_file_next[30][6] ), .D(\reg_file_next[31][6] ), .S0(n2236), .S1(
        n2219), .Y(n2719) );
  MXI4XL U2923 ( .A(\reg_file_next[12][7] ), .B(\reg_file_next[13][7] ), .C(
        \reg_file_next[14][7] ), .D(\reg_file_next[15][7] ), .S0(n2237), .S1(
        n2219), .Y(n2731) );
  MXI4XL U2924 ( .A(\reg_file_next[28][7] ), .B(\reg_file_next[29][7] ), .C(
        \reg_file_next[30][7] ), .D(\reg_file_next[31][7] ), .S0(n2237), .S1(
        n2219), .Y(n2727) );
  MXI4XL U2925 ( .A(\reg_file_next[12][8] ), .B(\reg_file_next[13][8] ), .C(
        \reg_file_next[14][8] ), .D(\reg_file_next[15][8] ), .S0(n2238), .S1(
        n2220), .Y(n2739) );
  MXI4XL U2926 ( .A(\reg_file_next[28][8] ), .B(\reg_file_next[29][8] ), .C(
        \reg_file_next[30][8] ), .D(\reg_file_next[31][8] ), .S0(n2237), .S1(
        n2219), .Y(n2735) );
  MXI4XL U2927 ( .A(\reg_file_next[12][9] ), .B(\reg_file_next[13][9] ), .C(
        \reg_file_next[14][9] ), .D(\reg_file_next[15][9] ), .S0(n2238), .S1(
        n2220), .Y(n2747) );
  MXI4XL U2928 ( .A(\reg_file_next[28][9] ), .B(\reg_file_next[29][9] ), .C(
        \reg_file_next[30][9] ), .D(\reg_file_next[31][9] ), .S0(n2238), .S1(
        n2220), .Y(n2743) );
  MXI4XL U2929 ( .A(\reg_file_next[12][10] ), .B(\reg_file_next[13][10] ), .C(
        \reg_file_next[14][10] ), .D(\reg_file_next[15][10] ), .S0(n2239), 
        .S1(n2220), .Y(n2755) );
  MXI4XL U2930 ( .A(\reg_file_next[28][10] ), .B(\reg_file_next[29][10] ), .C(
        \reg_file_next[30][10] ), .D(\reg_file_next[31][10] ), .S0(n2239), 
        .S1(n2220), .Y(n2751) );
  MXI4XL U2931 ( .A(\reg_file_next[12][11] ), .B(\reg_file_next[13][11] ), .C(
        \reg_file_next[14][11] ), .D(\reg_file_next[15][11] ), .S0(n2240), 
        .S1(n2221), .Y(n2763) );
  MXI4XL U2932 ( .A(\reg_file_next[28][11] ), .B(\reg_file_next[29][11] ), .C(
        \reg_file_next[30][11] ), .D(\reg_file_next[31][11] ), .S0(n2239), 
        .S1(n2221), .Y(n2759) );
  MXI4XL U2933 ( .A(\reg_file_next[12][12] ), .B(\reg_file_next[13][12] ), .C(
        \reg_file_next[14][12] ), .D(\reg_file_next[15][12] ), .S0(n2240), 
        .S1(n2221), .Y(n2771) );
  MXI4XL U2934 ( .A(\reg_file_next[28][12] ), .B(\reg_file_next[29][12] ), .C(
        \reg_file_next[30][12] ), .D(\reg_file_next[31][12] ), .S0(n2240), 
        .S1(n2221), .Y(n2767) );
  MXI4XL U2935 ( .A(\reg_file_next[12][13] ), .B(\reg_file_next[13][13] ), .C(
        \reg_file_next[14][13] ), .D(\reg_file_next[15][13] ), .S0(n2241), 
        .S1(n2222), .Y(n2779) );
  MXI4XL U2936 ( .A(\reg_file_next[28][13] ), .B(\reg_file_next[29][13] ), .C(
        \reg_file_next[30][13] ), .D(\reg_file_next[31][13] ), .S0(n2240), 
        .S1(n2221), .Y(n2775) );
  MXI4XL U2937 ( .A(\reg_file_next[12][14] ), .B(\reg_file_next[13][14] ), .C(
        \reg_file_next[14][14] ), .D(\reg_file_next[15][14] ), .S0(n2241), 
        .S1(n2222), .Y(n2787) );
  MXI4XL U2938 ( .A(\reg_file_next[28][14] ), .B(\reg_file_next[29][14] ), .C(
        \reg_file_next[30][14] ), .D(\reg_file_next[31][14] ), .S0(n2241), 
        .S1(n2222), .Y(n2783) );
  MXI4XL U2939 ( .A(\reg_file_next[12][15] ), .B(\reg_file_next[13][15] ), .C(
        \reg_file_next[14][15] ), .D(\reg_file_next[15][15] ), .S0(n2237), 
        .S1(n2222), .Y(n2795) );
  MXI4XL U2940 ( .A(\reg_file_next[28][15] ), .B(\reg_file_next[29][15] ), .C(
        \reg_file_next[30][15] ), .D(\reg_file_next[31][15] ), .S0(n2230), 
        .S1(n2222), .Y(n2791) );
  MXI4XL U2941 ( .A(\reg_file_next[12][16] ), .B(\reg_file_next[13][16] ), .C(
        \reg_file_next[14][16] ), .D(\reg_file_next[15][16] ), .S0(n2224), 
        .S1(n2210), .Y(n2803) );
  MXI4XL U2942 ( .A(\reg_file_next[28][16] ), .B(\reg_file_next[29][16] ), .C(
        \reg_file_next[30][16] ), .D(\reg_file_next[31][16] ), .S0(n2228), 
        .S1(n2213), .Y(n2799) );
  MXI4XL U2943 ( .A(\reg_file_next[12][17] ), .B(\reg_file_next[13][17] ), .C(
        \reg_file_next[14][17] ), .D(\reg_file_next[15][17] ), .S0(n2225), 
        .S1(n2210), .Y(n2811) );
  MXI4XL U2944 ( .A(\reg_file_next[28][17] ), .B(\reg_file_next[29][17] ), .C(
        \reg_file_next[30][17] ), .D(\reg_file_next[31][17] ), .S0(n2224), 
        .S1(n2210), .Y(n2807) );
  MXI4XL U2945 ( .A(\reg_file_next[12][18] ), .B(\reg_file_next[13][18] ), .C(
        \reg_file_next[14][18] ), .D(\reg_file_next[15][18] ), .S0(n2225), 
        .S1(n2211), .Y(n2819) );
  MXI4XL U2946 ( .A(\reg_file_next[28][18] ), .B(\reg_file_next[29][18] ), .C(
        \reg_file_next[30][18] ), .D(\reg_file_next[31][18] ), .S0(n2225), 
        .S1(n2211), .Y(n2815) );
  MXI4XL U2947 ( .A(\reg_file_next[12][19] ), .B(\reg_file_next[13][19] ), .C(
        \reg_file_next[14][19] ), .D(\reg_file_next[15][19] ), .S0(n2226), 
        .S1(n2211), .Y(n2827) );
  MXI4XL U2948 ( .A(\reg_file_next[28][19] ), .B(\reg_file_next[29][19] ), .C(
        \reg_file_next[30][19] ), .D(\reg_file_next[31][19] ), .S0(n2226), 
        .S1(n2211), .Y(n2823) );
  MXI4XL U2949 ( .A(\reg_file_next[12][20] ), .B(\reg_file_next[13][20] ), .C(
        \reg_file_next[14][20] ), .D(\reg_file_next[15][20] ), .S0(n2226), 
        .S1(n2212), .Y(n2835) );
  MXI4XL U2950 ( .A(\reg_file_next[28][20] ), .B(\reg_file_next[29][20] ), .C(
        \reg_file_next[30][20] ), .D(\reg_file_next[31][20] ), .S0(n2226), 
        .S1(n2211), .Y(n2831) );
  MXI4XL U2951 ( .A(\reg_file_next[12][21] ), .B(\reg_file_next[13][21] ), .C(
        \reg_file_next[14][21] ), .D(\reg_file_next[15][21] ), .S0(n2227), 
        .S1(n2212), .Y(n2843) );
  MXI4XL U2952 ( .A(\reg_file_next[28][21] ), .B(\reg_file_next[29][21] ), .C(
        \reg_file_next[30][21] ), .D(\reg_file_next[31][21] ), .S0(n2227), 
        .S1(n2212), .Y(n2839) );
  MXI4XL U2953 ( .A(\reg_file_next[12][22] ), .B(\reg_file_next[13][22] ), .C(
        \reg_file_next[14][22] ), .D(\reg_file_next[15][22] ), .S0(n2228), 
        .S1(n2212), .Y(n2851) );
  MXI4XL U2954 ( .A(\reg_file_next[28][22] ), .B(\reg_file_next[29][22] ), .C(
        \reg_file_next[30][22] ), .D(\reg_file_next[31][22] ), .S0(n2227), 
        .S1(n2212), .Y(n2847) );
  MXI4XL U2955 ( .A(\reg_file_next[12][23] ), .B(\reg_file_next[13][23] ), .C(
        \reg_file_next[14][23] ), .D(\reg_file_next[15][23] ), .S0(n2228), 
        .S1(n2213), .Y(n2859) );
  MXI4XL U2956 ( .A(\reg_file_next[28][23] ), .B(\reg_file_next[29][23] ), .C(
        \reg_file_next[30][23] ), .D(\reg_file_next[31][23] ), .S0(n2228), 
        .S1(n2213), .Y(n2855) );
  MXI4XL U2957 ( .A(\reg_file_next[12][24] ), .B(\reg_file_next[13][24] ), .C(
        \reg_file_next[14][24] ), .D(\reg_file_next[15][24] ), .S0(n2229), 
        .S1(n2213), .Y(n2867) );
  MXI4XL U2958 ( .A(\reg_file_next[28][24] ), .B(\reg_file_next[29][24] ), .C(
        \reg_file_next[30][24] ), .D(\reg_file_next[31][24] ), .S0(n2233), 
        .S1(n2216), .Y(n2863) );
  MXI4XL U2959 ( .A(\reg_file_next[12][25] ), .B(\reg_file_next[13][25] ), .C(
        \reg_file_next[14][25] ), .D(\reg_file_next[15][25] ), .S0(n2229), 
        .S1(n2214), .Y(n2875) );
  MXI4XL U2960 ( .A(\reg_file_next[28][25] ), .B(\reg_file_next[29][25] ), .C(
        \reg_file_next[30][25] ), .D(\reg_file_next[31][25] ), .S0(n2229), 
        .S1(n2213), .Y(n2871) );
  MXI4XL U2961 ( .A(\reg_file_next[12][26] ), .B(\reg_file_next[13][26] ), .C(
        \reg_file_next[14][26] ), .D(\reg_file_next[15][26] ), .S0(n2230), 
        .S1(n2214), .Y(n2883) );
  MXI4XL U2962 ( .A(\reg_file_next[28][26] ), .B(\reg_file_next[29][26] ), .C(
        \reg_file_next[30][26] ), .D(\reg_file_next[31][26] ), .S0(n2230), 
        .S1(n2214), .Y(n2879) );
  MXI4XL U2963 ( .A(\reg_file_next[12][27] ), .B(\reg_file_next[13][27] ), .C(
        \reg_file_next[14][27] ), .D(\reg_file_next[15][27] ), .S0(n2230), 
        .S1(n2214), .Y(n2891) );
  MXI4XL U2964 ( .A(\reg_file_next[28][27] ), .B(\reg_file_next[29][27] ), .C(
        \reg_file_next[30][27] ), .D(\reg_file_next[31][27] ), .S0(n2230), 
        .S1(n2214), .Y(n2887) );
  MXI4XL U2965 ( .A(\reg_file_next[12][28] ), .B(\reg_file_next[13][28] ), .C(
        \reg_file_next[14][28] ), .D(\reg_file_next[15][28] ), .S0(n2231), 
        .S1(n2215), .Y(n2899) );
  MXI4XL U2966 ( .A(\reg_file_next[28][28] ), .B(\reg_file_next[29][28] ), .C(
        \reg_file_next[30][28] ), .D(\reg_file_next[31][28] ), .S0(n2231), 
        .S1(n2215), .Y(n2895) );
  MXI4XL U2967 ( .A(\reg_file_next[12][29] ), .B(\reg_file_next[13][29] ), .C(
        \reg_file_next[14][29] ), .D(\reg_file_next[15][29] ), .S0(n2232), 
        .S1(n2215), .Y(n2907) );
  MXI4XL U2968 ( .A(\reg_file_next[28][29] ), .B(\reg_file_next[29][29] ), .C(
        \reg_file_next[30][29] ), .D(\reg_file_next[31][29] ), .S0(n2231), 
        .S1(n2215), .Y(n2903) );
  MXI4XL U2969 ( .A(\reg_file_next[12][30] ), .B(\reg_file_next[13][30] ), .C(
        \reg_file_next[14][30] ), .D(\reg_file_next[15][30] ), .S0(n2232), 
        .S1(n2216), .Y(n2915) );
  MXI4XL U2970 ( .A(\reg_file_next[28][30] ), .B(\reg_file_next[29][30] ), .C(
        \reg_file_next[30][30] ), .D(\reg_file_next[31][30] ), .S0(n2232), 
        .S1(n2215), .Y(n2911) );
  MXI4XL U2971 ( .A(\reg_file_next[12][31] ), .B(\reg_file_next[13][31] ), .C(
        \reg_file_next[14][31] ), .D(\reg_file_next[15][31] ), .S0(n2233), 
        .S1(n2216), .Y(n2923) );
  MXI4XL U2972 ( .A(\reg_file_next[28][31] ), .B(\reg_file_next[29][31] ), .C(
        \reg_file_next[30][31] ), .D(\reg_file_next[31][31] ), .S0(n2232), 
        .S1(n2216), .Y(n2919) );
  MXI4XL U2973 ( .A(\reg_file_next[12][0] ), .B(\reg_file_next[13][0] ), .C(
        \reg_file_next[14][0] ), .D(\reg_file_next[15][0] ), .S0(n2262), .S1(
        n2243), .Y(n2355) );
  MXI4XL U2974 ( .A(\reg_file_next[28][0] ), .B(\reg_file_next[29][0] ), .C(
        \reg_file_next[30][0] ), .D(\reg_file_next[31][0] ), .S0(n2253), .S1(
        n2242), .Y(n2351) );
  MXI4XL U2975 ( .A(\reg_file_next[12][1] ), .B(\reg_file_next[13][1] ), .C(
        \reg_file_next[14][1] ), .D(\reg_file_next[15][1] ), .S0(n2263), .S1(
        n2252), .Y(n2363) );
  MXI4XL U2976 ( .A(\reg_file_next[28][1] ), .B(\reg_file_next[29][1] ), .C(
        \reg_file_next[30][1] ), .D(\reg_file_next[31][1] ), .S0(n2262), .S1(
        n2247), .Y(n2359) );
  MXI4XL U2977 ( .A(\reg_file_next[12][2] ), .B(\reg_file_next[13][2] ), .C(
        \reg_file_next[14][2] ), .D(\reg_file_next[15][2] ), .S0(n2263), .S1(
        n2247), .Y(n2371) );
  MXI4XL U2978 ( .A(\reg_file_next[28][2] ), .B(\reg_file_next[29][2] ), .C(
        \reg_file_next[30][2] ), .D(\reg_file_next[31][2] ), .S0(n2263), .S1(
        n2247), .Y(n2367) );
  MXI4XL U2979 ( .A(\reg_file_next[12][3] ), .B(\reg_file_next[13][3] ), .C(
        \reg_file_next[14][3] ), .D(\reg_file_next[15][3] ), .S0(n2264), .S1(
        n2247), .Y(n2379) );
  MXI4XL U2980 ( .A(\reg_file_next[28][3] ), .B(\reg_file_next[29][3] ), .C(
        \reg_file_next[30][3] ), .D(\reg_file_next[31][3] ), .S0(n2264), .S1(
        n2247), .Y(n2375) );
  MXI4XL U2981 ( .A(\reg_file_next[12][4] ), .B(\reg_file_next[13][4] ), .C(
        \reg_file_next[14][4] ), .D(\reg_file_next[15][4] ), .S0(n2264), .S1(
        n2248), .Y(n2387) );
  MXI4XL U2982 ( .A(\reg_file_next[28][4] ), .B(\reg_file_next[29][4] ), .C(
        \reg_file_next[30][4] ), .D(\reg_file_next[31][4] ), .S0(n2264), .S1(
        n2247), .Y(n2383) );
  MXI4XL U2983 ( .A(\reg_file_next[12][5] ), .B(\reg_file_next[13][5] ), .C(
        \reg_file_next[14][5] ), .D(\reg_file_next[15][5] ), .S0(n2265), .S1(
        n2248), .Y(n2395) );
  MXI4XL U2984 ( .A(\reg_file_next[28][5] ), .B(\reg_file_next[29][5] ), .C(
        \reg_file_next[30][5] ), .D(\reg_file_next[31][5] ), .S0(n2265), .S1(
        n2248), .Y(n2391) );
  MXI4XL U2985 ( .A(\reg_file_next[12][6] ), .B(\reg_file_next[13][6] ), .C(
        \reg_file_next[14][6] ), .D(\reg_file_next[15][6] ), .S0(n2266), .S1(
        n2248), .Y(n2403) );
  MXI4XL U2986 ( .A(\reg_file_next[28][6] ), .B(\reg_file_next[29][6] ), .C(
        \reg_file_next[30][6] ), .D(\reg_file_next[31][6] ), .S0(n2265), .S1(
        n2248), .Y(n2399) );
  MXI4XL U2987 ( .A(\reg_file_next[12][7] ), .B(\reg_file_next[13][7] ), .C(
        \reg_file_next[14][7] ), .D(\reg_file_next[15][7] ), .S0(n2266), .S1(
        n2249), .Y(n2411) );
  MXI4XL U2988 ( .A(\reg_file_next[28][7] ), .B(\reg_file_next[29][7] ), .C(
        \reg_file_next[30][7] ), .D(\reg_file_next[31][7] ), .S0(n2266), .S1(
        n2249), .Y(n2407) );
  MXI4XL U2989 ( .A(\reg_file_next[12][8] ), .B(\reg_file_next[13][8] ), .C(
        \reg_file_next[14][8] ), .D(\reg_file_next[15][8] ), .S0(n2267), .S1(
        n2249), .Y(n2419) );
  MXI4XL U2990 ( .A(\reg_file_next[28][8] ), .B(\reg_file_next[29][8] ), .C(
        \reg_file_next[30][8] ), .D(\reg_file_next[31][8] ), .S0(n2266), .S1(
        n2249), .Y(n2415) );
  MXI4XL U2991 ( .A(\reg_file_next[12][9] ), .B(\reg_file_next[13][9] ), .C(
        \reg_file_next[14][9] ), .D(\reg_file_next[15][9] ), .S0(n2267), .S1(
        n2250), .Y(n2427) );
  MXI4XL U2992 ( .A(\reg_file_next[28][9] ), .B(\reg_file_next[29][9] ), .C(
        \reg_file_next[30][9] ), .D(\reg_file_next[31][9] ), .S0(n2267), .S1(
        n2249), .Y(n2423) );
  MXI4XL U2993 ( .A(\reg_file_next[12][10] ), .B(\reg_file_next[13][10] ), .C(
        \reg_file_next[14][10] ), .D(\reg_file_next[15][10] ), .S0(n2268), 
        .S1(n2250), .Y(n2435) );
  MXI4XL U2994 ( .A(\reg_file_next[28][10] ), .B(\reg_file_next[29][10] ), .C(
        \reg_file_next[30][10] ), .D(\reg_file_next[31][10] ), .S0(n2268), 
        .S1(n2250), .Y(n2431) );
  MXI4XL U2995 ( .A(\reg_file_next[12][11] ), .B(\reg_file_next[13][11] ), .C(
        \reg_file_next[14][11] ), .D(\reg_file_next[15][11] ), .S0(n2269), 
        .S1(n2250), .Y(n2443) );
  MXI4XL U2996 ( .A(\reg_file_next[28][11] ), .B(\reg_file_next[29][11] ), .C(
        \reg_file_next[30][11] ), .D(\reg_file_next[31][11] ), .S0(n2268), 
        .S1(n2250), .Y(n2439) );
  MXI4XL U2997 ( .A(\reg_file_next[12][12] ), .B(\reg_file_next[13][12] ), .C(
        \reg_file_next[14][12] ), .D(\reg_file_next[15][12] ), .S0(n2269), 
        .S1(n2251), .Y(n2451) );
  MXI4XL U2998 ( .A(\reg_file_next[28][12] ), .B(\reg_file_next[29][12] ), .C(
        \reg_file_next[30][12] ), .D(\reg_file_next[31][12] ), .S0(n2269), 
        .S1(n2251), .Y(n2447) );
  MXI4XL U2999 ( .A(\reg_file_next[12][13] ), .B(\reg_file_next[13][13] ), .C(
        \reg_file_next[14][13] ), .D(\reg_file_next[15][13] ), .S0(n2270), 
        .S1(n2251), .Y(n2459) );
  MXI4XL U3000 ( .A(\reg_file_next[28][13] ), .B(\reg_file_next[29][13] ), .C(
        \reg_file_next[30][13] ), .D(\reg_file_next[31][13] ), .S0(n2269), 
        .S1(n2251), .Y(n2455) );
  MXI4XL U3001 ( .A(\reg_file_next[12][14] ), .B(\reg_file_next[13][14] ), .C(
        \reg_file_next[14][14] ), .D(\reg_file_next[15][14] ), .S0(n2270), 
        .S1(n2251), .Y(n2467) );
  MXI4XL U3002 ( .A(\reg_file_next[28][14] ), .B(\reg_file_next[29][14] ), .C(
        \reg_file_next[30][14] ), .D(\reg_file_next[31][14] ), .S0(n2270), 
        .S1(n2251), .Y(n2463) );
  MXI4XL U3003 ( .A(\reg_file_next[12][15] ), .B(\reg_file_next[13][15] ), .C(
        \reg_file_next[14][15] ), .D(\reg_file_next[15][15] ), .S0(n2257), 
        .S1(n2252), .Y(n2475) );
  MXI4XL U3004 ( .A(\reg_file_next[28][15] ), .B(\reg_file_next[29][15] ), .C(
        \reg_file_next[30][15] ), .D(\reg_file_next[31][15] ), .S0(n2260), 
        .S1(n2252), .Y(n2471) );
  MXI4XL U3005 ( .A(\reg_file_next[12][16] ), .B(\reg_file_next[13][16] ), .C(
        \reg_file_next[14][16] ), .D(\reg_file_next[15][16] ), .S0(n2253), 
        .S1(n2242), .Y(n2483) );
  MXI4XL U3006 ( .A(\reg_file_next[28][16] ), .B(\reg_file_next[29][16] ), .C(
        \reg_file_next[30][16] ), .D(\reg_file_next[31][16] ), .S0(n2257), 
        .S1(n2244), .Y(n2479) );
  MXI4XL U3007 ( .A(\reg_file_next[12][17] ), .B(\reg_file_next[13][17] ), .C(
        \reg_file_next[14][17] ), .D(\reg_file_next[15][17] ), .S0(n2254), 
        .S1(n2242), .Y(n2491) );
  MXI4XL U3008 ( .A(\reg_file_next[28][17] ), .B(\reg_file_next[29][17] ), .C(
        \reg_file_next[30][17] ), .D(\reg_file_next[31][17] ), .S0(n2253), 
        .S1(n2242), .Y(n2487) );
  MXI4XL U3009 ( .A(\reg_file_next[12][18] ), .B(\reg_file_next[13][18] ), .C(
        \reg_file_next[14][18] ), .D(\reg_file_next[15][18] ), .S0(n2254), 
        .S1(n2243), .Y(n2499) );
  MXI4XL U3010 ( .A(\reg_file_next[28][18] ), .B(\reg_file_next[29][18] ), .C(
        \reg_file_next[30][18] ), .D(\reg_file_next[31][18] ), .S0(n2254), 
        .S1(n2243), .Y(n2495) );
  MXI4XL U3011 ( .A(\reg_file_next[12][19] ), .B(\reg_file_next[13][19] ), .C(
        \reg_file_next[14][19] ), .D(\reg_file_next[15][19] ), .S0(n2255), 
        .S1(n2243), .Y(n2507) );
  MXI4XL U3012 ( .A(\reg_file_next[28][19] ), .B(\reg_file_next[29][19] ), .C(
        \reg_file_next[30][19] ), .D(\reg_file_next[31][19] ), .S0(n2255), 
        .S1(n2243), .Y(n2503) );
  MXI4XL U3013 ( .A(\reg_file_next[12][20] ), .B(\reg_file_next[13][20] ), .C(
        \reg_file_next[14][20] ), .D(\reg_file_next[15][20] ), .S0(n2255), 
        .S1(n2247), .Y(n2515) );
  MXI4XL U3014 ( .A(\reg_file_next[28][20] ), .B(\reg_file_next[29][20] ), .C(
        \reg_file_next[30][20] ), .D(\reg_file_next[31][20] ), .S0(n2255), 
        .S1(n2243), .Y(n2511) );
  MXI4XL U3015 ( .A(\reg_file_next[12][21] ), .B(\reg_file_next[13][21] ), .C(
        \reg_file_next[14][21] ), .D(\reg_file_next[15][21] ), .S0(n2256), 
        .S1(n2245), .Y(n2523) );
  MXI4XL U3016 ( .A(\reg_file_next[28][21] ), .B(\reg_file_next[29][21] ), .C(
        \reg_file_next[30][21] ), .D(\reg_file_next[31][21] ), .S0(n2256), 
        .S1(n2249), .Y(n2519) );
  MXI4XL U3017 ( .A(\reg_file_next[12][22] ), .B(\reg_file_next[13][22] ), .C(
        \reg_file_next[14][22] ), .D(\reg_file_next[15][22] ), .S0(n2257), 
        .S1(n2246), .Y(n2531) );
  MXI4XL U3018 ( .A(\reg_file_next[28][22] ), .B(\reg_file_next[29][22] ), .C(
        \reg_file_next[30][22] ), .D(\reg_file_next[31][22] ), .S0(n2256), 
        .S1(n2244), .Y(n2527) );
  MXI4XL U3019 ( .A(\reg_file_next[12][23] ), .B(\reg_file_next[13][23] ), .C(
        \reg_file_next[14][23] ), .D(\reg_file_next[15][23] ), .S0(n2257), 
        .S1(n2244), .Y(n2539) );
  MXI4XL U3020 ( .A(\reg_file_next[28][23] ), .B(\reg_file_next[29][23] ), .C(
        \reg_file_next[30][23] ), .D(\reg_file_next[31][23] ), .S0(n2257), 
        .S1(n2244), .Y(n2535) );
  MXI4XL U3021 ( .A(\reg_file_next[12][24] ), .B(\reg_file_next[13][24] ), .C(
        \reg_file_next[14][24] ), .D(\reg_file_next[15][24] ), .S0(n2258), 
        .S1(n2244), .Y(n2547) );
  MXI4XL U3022 ( .A(\reg_file_next[28][24] ), .B(\reg_file_next[29][24] ), .C(
        \reg_file_next[30][24] ), .D(\reg_file_next[31][24] ), .S0(n2262), 
        .S1(n2245), .Y(n2543) );
  MXI4XL U3023 ( .A(\reg_file_next[12][25] ), .B(\reg_file_next[13][25] ), .C(
        \reg_file_next[14][25] ), .D(\reg_file_next[15][25] ), .S0(n2258), 
        .S1(n2244), .Y(n2555) );
  MXI4XL U3024 ( .A(\reg_file_next[28][25] ), .B(\reg_file_next[29][25] ), .C(
        \reg_file_next[30][25] ), .D(\reg_file_next[31][25] ), .S0(n2258), 
        .S1(n2244), .Y(n2551) );
  MXI4XL U3025 ( .A(\reg_file_next[12][26] ), .B(\reg_file_next[13][26] ), .C(
        \reg_file_next[14][26] ), .D(\reg_file_next[15][26] ), .S0(n2259), 
        .S1(n2245), .Y(n2563) );
  MXI4XL U3026 ( .A(\reg_file_next[28][26] ), .B(\reg_file_next[29][26] ), .C(
        \reg_file_next[30][26] ), .D(\reg_file_next[31][26] ), .S0(n2259), 
        .S1(n2245), .Y(n2559) );
  MXI4XL U3027 ( .A(\reg_file_next[12][27] ), .B(\reg_file_next[13][27] ), .C(
        \reg_file_next[14][27] ), .D(\reg_file_next[15][27] ), .S0(n2259), 
        .S1(n2245), .Y(n2571) );
  MXI4XL U3028 ( .A(\reg_file_next[28][27] ), .B(\reg_file_next[29][27] ), .C(
        \reg_file_next[30][27] ), .D(\reg_file_next[31][27] ), .S0(n2259), 
        .S1(n2245), .Y(n2567) );
  MXI4XL U3029 ( .A(\reg_file_next[12][28] ), .B(\reg_file_next[13][28] ), .C(
        \reg_file_next[14][28] ), .D(\reg_file_next[15][28] ), .S0(n2260), 
        .S1(n2246), .Y(n2579) );
  MXI4XL U3030 ( .A(\reg_file_next[28][28] ), .B(\reg_file_next[29][28] ), .C(
        \reg_file_next[30][28] ), .D(\reg_file_next[31][28] ), .S0(n2260), 
        .S1(n2245), .Y(n2575) );
  MXI4XL U3031 ( .A(\reg_file_next[12][29] ), .B(\reg_file_next[13][29] ), .C(
        \reg_file_next[14][29] ), .D(\reg_file_next[15][29] ), .S0(n2261), 
        .S1(n2246), .Y(n2587) );
  MXI4XL U3032 ( .A(\reg_file_next[28][29] ), .B(\reg_file_next[29][29] ), .C(
        \reg_file_next[30][29] ), .D(\reg_file_next[31][29] ), .S0(n2260), 
        .S1(n2246), .Y(n2583) );
  MXI4XL U3033 ( .A(\reg_file_next[12][30] ), .B(\reg_file_next[13][30] ), .C(
        \reg_file_next[14][30] ), .D(\reg_file_next[15][30] ), .S0(n2261), 
        .S1(n2246), .Y(n2595) );
  MXI4XL U3034 ( .A(\reg_file_next[28][30] ), .B(\reg_file_next[29][30] ), .C(
        \reg_file_next[30][30] ), .D(\reg_file_next[31][30] ), .S0(n2261), 
        .S1(n2246), .Y(n2591) );
  MXI4XL U3035 ( .A(\reg_file_next[12][31] ), .B(\reg_file_next[13][31] ), .C(
        \reg_file_next[14][31] ), .D(\reg_file_next[15][31] ), .S0(n2262), 
        .S1(n2249), .Y(n2603) );
  MXI4XL U3036 ( .A(\reg_file_next[28][31] ), .B(\reg_file_next[29][31] ), .C(
        \reg_file_next[30][31] ), .D(\reg_file_next[31][31] ), .S0(n2261), 
        .S1(n2246), .Y(n2599) );
  MXI4XL U3037 ( .A(\reg_file_next[8][0] ), .B(\reg_file_next[9][0] ), .C(
        \reg_file_next[10][0] ), .D(\reg_file_next[11][0] ), .S0(n2233), .S1(
        n2216), .Y(n2676) );
  MXI4XL U3038 ( .A(\reg_file_next[8][1] ), .B(\reg_file_next[9][1] ), .C(
        \reg_file_next[10][1] ), .D(\reg_file_next[11][1] ), .S0(n2234), .S1(
        n2217), .Y(n2684) );
  MXI4XL U3039 ( .A(\reg_file_next[8][2] ), .B(\reg_file_next[9][2] ), .C(
        \reg_file_next[10][2] ), .D(\reg_file_next[11][2] ), .S0(n2234), .S1(
        n2217), .Y(n2692) );
  MXI4XL U3040 ( .A(\reg_file_next[8][3] ), .B(\reg_file_next[9][3] ), .C(
        \reg_file_next[10][3] ), .D(\reg_file_next[11][3] ), .S0(n2235), .S1(
        n2218), .Y(n2700) );
  MXI4XL U3041 ( .A(\reg_file_next[8][4] ), .B(\reg_file_next[9][4] ), .C(
        \reg_file_next[10][4] ), .D(\reg_file_next[11][4] ), .S0(n2236), .S1(
        n2218), .Y(n2708) );
  MXI4XL U3042 ( .A(\reg_file_next[8][5] ), .B(\reg_file_next[9][5] ), .C(
        \reg_file_next[10][5] ), .D(\reg_file_next[11][5] ), .S0(n2236), .S1(
        n2218), .Y(n2716) );
  MXI4XL U3043 ( .A(\reg_file_next[8][6] ), .B(\reg_file_next[9][6] ), .C(
        \reg_file_next[10][6] ), .D(\reg_file_next[11][6] ), .S0(n2237), .S1(
        n2219), .Y(n2724) );
  MXI4XL U3044 ( .A(\reg_file_next[8][7] ), .B(\reg_file_next[9][7] ), .C(
        \reg_file_next[10][7] ), .D(\reg_file_next[11][7] ), .S0(n2237), .S1(
        n2219), .Y(n2732) );
  MXI4XL U3045 ( .A(\reg_file_next[8][8] ), .B(\reg_file_next[9][8] ), .C(
        \reg_file_next[10][8] ), .D(\reg_file_next[11][8] ), .S0(n2238), .S1(
        n2220), .Y(n2740) );
  MXI4XL U3046 ( .A(\reg_file_next[8][9] ), .B(\reg_file_next[9][9] ), .C(
        \reg_file_next[10][9] ), .D(\reg_file_next[11][9] ), .S0(n2238), .S1(
        n2220), .Y(n2748) );
  MXI4XL U3047 ( .A(\reg_file_next[8][10] ), .B(\reg_file_next[9][10] ), .C(
        \reg_file_next[10][10] ), .D(\reg_file_next[11][10] ), .S0(n2239), 
        .S1(n2220), .Y(n2756) );
  MXI4XL U3048 ( .A(\reg_file_next[8][11] ), .B(\reg_file_next[9][11] ), .C(
        \reg_file_next[10][11] ), .D(\reg_file_next[11][11] ), .S0(n2240), 
        .S1(n2221), .Y(n2764) );
  MXI4XL U3049 ( .A(\reg_file_next[8][12] ), .B(\reg_file_next[9][12] ), .C(
        \reg_file_next[10][12] ), .D(\reg_file_next[11][12] ), .S0(n2240), 
        .S1(n2221), .Y(n2772) );
  MXI4XL U3050 ( .A(\reg_file_next[8][13] ), .B(\reg_file_next[9][13] ), .C(
        \reg_file_next[10][13] ), .D(\reg_file_next[11][13] ), .S0(n2241), 
        .S1(n2222), .Y(n2780) );
  MXI4XL U3051 ( .A(\reg_file_next[8][14] ), .B(\reg_file_next[9][14] ), .C(
        \reg_file_next[10][14] ), .D(\reg_file_next[11][14] ), .S0(n2241), 
        .S1(n2222), .Y(n2788) );
  MXI4XL U3052 ( .A(\reg_file_next[8][15] ), .B(\reg_file_next[9][15] ), .C(
        \reg_file_next[10][15] ), .D(\reg_file_next[11][15] ), .S0(n2231), 
        .S1(n2222), .Y(n2796) );
  MXI4XL U3053 ( .A(\reg_file_next[8][16] ), .B(\reg_file_next[9][16] ), .C(
        \reg_file_next[10][16] ), .D(\reg_file_next[11][16] ), .S0(n2224), 
        .S1(n2210), .Y(n2804) );
  MXI4XL U3054 ( .A(\reg_file_next[8][17] ), .B(\reg_file_next[9][17] ), .C(
        \reg_file_next[10][17] ), .D(\reg_file_next[11][17] ), .S0(n2225), 
        .S1(n2210), .Y(n2812) );
  MXI4XL U3055 ( .A(\reg_file_next[8][18] ), .B(\reg_file_next[9][18] ), .C(
        \reg_file_next[10][18] ), .D(\reg_file_next[11][18] ), .S0(n2225), 
        .S1(n2211), .Y(n2820) );
  MXI4XL U3056 ( .A(\reg_file_next[8][19] ), .B(\reg_file_next[9][19] ), .C(
        \reg_file_next[10][19] ), .D(\reg_file_next[11][19] ), .S0(n2226), 
        .S1(n2211), .Y(n2828) );
  MXI4XL U3057 ( .A(\reg_file_next[8][20] ), .B(\reg_file_next[9][20] ), .C(
        \reg_file_next[10][20] ), .D(\reg_file_next[11][20] ), .S0(n2226), 
        .S1(n2212), .Y(n2836) );
  MXI4XL U3058 ( .A(\reg_file_next[8][21] ), .B(\reg_file_next[9][21] ), .C(
        \reg_file_next[10][21] ), .D(\reg_file_next[11][21] ), .S0(n2227), 
        .S1(n2212), .Y(n2844) );
  MXI4XL U3059 ( .A(\reg_file_next[8][22] ), .B(\reg_file_next[9][22] ), .C(
        \reg_file_next[10][22] ), .D(\reg_file_next[11][22] ), .S0(n2228), 
        .S1(n2212), .Y(n2852) );
  MXI4XL U3060 ( .A(\reg_file_next[8][23] ), .B(\reg_file_next[9][23] ), .C(
        \reg_file_next[10][23] ), .D(\reg_file_next[11][23] ), .S0(n2228), 
        .S1(n2213), .Y(n2860) );
  MXI4XL U3061 ( .A(\reg_file_next[8][24] ), .B(\reg_file_next[9][24] ), .C(
        \reg_file_next[10][24] ), .D(\reg_file_next[11][24] ), .S0(n2229), 
        .S1(n2213), .Y(n2868) );
  MXI4XL U3062 ( .A(\reg_file_next[8][25] ), .B(\reg_file_next[9][25] ), .C(
        \reg_file_next[10][25] ), .D(\reg_file_next[11][25] ), .S0(n2229), 
        .S1(n2214), .Y(n2876) );
  MXI4XL U3063 ( .A(\reg_file_next[8][26] ), .B(\reg_file_next[9][26] ), .C(
        \reg_file_next[10][26] ), .D(\reg_file_next[11][26] ), .S0(n2230), 
        .S1(n2214), .Y(n2884) );
  MXI4XL U3064 ( .A(\reg_file_next[8][27] ), .B(\reg_file_next[9][27] ), .C(
        \reg_file_next[10][27] ), .D(\reg_file_next[11][27] ), .S0(n2230), 
        .S1(n2214), .Y(n2892) );
  MXI4XL U3065 ( .A(\reg_file_next[8][28] ), .B(\reg_file_next[9][28] ), .C(
        \reg_file_next[10][28] ), .D(\reg_file_next[11][28] ), .S0(n2231), 
        .S1(n2215), .Y(n2900) );
  MXI4XL U3066 ( .A(\reg_file_next[8][29] ), .B(\reg_file_next[9][29] ), .C(
        \reg_file_next[10][29] ), .D(\reg_file_next[11][29] ), .S0(n2232), 
        .S1(n2215), .Y(n2908) );
  MXI4XL U3067 ( .A(\reg_file_next[8][30] ), .B(\reg_file_next[9][30] ), .C(
        \reg_file_next[10][30] ), .D(\reg_file_next[11][30] ), .S0(n2232), 
        .S1(n2216), .Y(n2916) );
  MXI4XL U3068 ( .A(\reg_file_next[8][31] ), .B(\reg_file_next[9][31] ), .C(
        \reg_file_next[10][31] ), .D(\reg_file_next[11][31] ), .S0(n2233), 
        .S1(n2216), .Y(n2924) );
  MXI4XL U3069 ( .A(\reg_file_next[8][0] ), .B(\reg_file_next[9][0] ), .C(
        \reg_file_next[10][0] ), .D(\reg_file_next[11][0] ), .S0(n2262), .S1(
        n2244), .Y(n2356) );
  MXI4XL U3070 ( .A(\reg_file_next[8][1] ), .B(\reg_file_next[9][1] ), .C(
        \reg_file_next[10][1] ), .D(\reg_file_next[11][1] ), .S0(n2263), .S1(
        n2247), .Y(n2364) );
  MXI4XL U3071 ( .A(\reg_file_next[8][2] ), .B(\reg_file_next[9][2] ), .C(
        \reg_file_next[10][2] ), .D(\reg_file_next[11][2] ), .S0(n2263), .S1(
        n2247), .Y(n2372) );
  MXI4XL U3072 ( .A(\reg_file_next[8][3] ), .B(\reg_file_next[9][3] ), .C(
        \reg_file_next[10][3] ), .D(\reg_file_next[11][3] ), .S0(n2264), .S1(
        n2247), .Y(n2380) );
  MXI4XL U3073 ( .A(\reg_file_next[8][4] ), .B(\reg_file_next[9][4] ), .C(
        \reg_file_next[10][4] ), .D(\reg_file_next[11][4] ), .S0(n2265), .S1(
        n2248), .Y(n2388) );
  MXI4XL U3074 ( .A(\reg_file_next[8][5] ), .B(\reg_file_next[9][5] ), .C(
        \reg_file_next[10][5] ), .D(\reg_file_next[11][5] ), .S0(n2265), .S1(
        n2248), .Y(n2396) );
  MXI4XL U3075 ( .A(\reg_file_next[8][6] ), .B(\reg_file_next[9][6] ), .C(
        \reg_file_next[10][6] ), .D(\reg_file_next[11][6] ), .S0(n2266), .S1(
        n2248), .Y(n2404) );
  MXI4XL U3076 ( .A(\reg_file_next[8][7] ), .B(\reg_file_next[9][7] ), .C(
        \reg_file_next[10][7] ), .D(\reg_file_next[11][7] ), .S0(n2266), .S1(
        n2249), .Y(n2412) );
  MXI4XL U3077 ( .A(\reg_file_next[8][8] ), .B(\reg_file_next[9][8] ), .C(
        \reg_file_next[10][8] ), .D(\reg_file_next[11][8] ), .S0(n2267), .S1(
        n2249), .Y(n2420) );
  MXI4XL U3078 ( .A(\reg_file_next[8][9] ), .B(\reg_file_next[9][9] ), .C(
        \reg_file_next[10][9] ), .D(\reg_file_next[11][9] ), .S0(n2267), .S1(
        n2250), .Y(n2428) );
  MXI4XL U3079 ( .A(\reg_file_next[8][10] ), .B(\reg_file_next[9][10] ), .C(
        \reg_file_next[10][10] ), .D(\reg_file_next[11][10] ), .S0(n2268), 
        .S1(n2250), .Y(n2436) );
  MXI4XL U3080 ( .A(\reg_file_next[8][11] ), .B(\reg_file_next[9][11] ), .C(
        \reg_file_next[10][11] ), .D(\reg_file_next[11][11] ), .S0(n2269), 
        .S1(n2250), .Y(n2444) );
  MXI4XL U3081 ( .A(\reg_file_next[8][12] ), .B(\reg_file_next[9][12] ), .C(
        \reg_file_next[10][12] ), .D(\reg_file_next[11][12] ), .S0(n2269), 
        .S1(n2251), .Y(n2452) );
  MXI4XL U3082 ( .A(\reg_file_next[8][13] ), .B(\reg_file_next[9][13] ), .C(
        \reg_file_next[10][13] ), .D(\reg_file_next[11][13] ), .S0(n2270), 
        .S1(n2251), .Y(n2460) );
  MXI4XL U3083 ( .A(\reg_file_next[8][14] ), .B(\reg_file_next[9][14] ), .C(
        \reg_file_next[10][14] ), .D(\reg_file_next[11][14] ), .S0(n2270), 
        .S1(n2252), .Y(n2468) );
  MXI4XL U3084 ( .A(\reg_file_next[8][15] ), .B(\reg_file_next[9][15] ), .C(
        \reg_file_next[10][15] ), .D(\reg_file_next[11][15] ), .S0(n2258), 
        .S1(n2252), .Y(n2476) );
  MXI4XL U3085 ( .A(\reg_file_next[8][16] ), .B(\reg_file_next[9][16] ), .C(
        \reg_file_next[10][16] ), .D(\reg_file_next[11][16] ), .S0(n2253), 
        .S1(n2242), .Y(n2484) );
  MXI4XL U3086 ( .A(\reg_file_next[8][17] ), .B(\reg_file_next[9][17] ), .C(
        \reg_file_next[10][17] ), .D(\reg_file_next[11][17] ), .S0(n2254), 
        .S1(n2242), .Y(n2492) );
  MXI4XL U3087 ( .A(\reg_file_next[8][18] ), .B(\reg_file_next[9][18] ), .C(
        \reg_file_next[10][18] ), .D(\reg_file_next[11][18] ), .S0(n2254), 
        .S1(n2243), .Y(n2500) );
  MXI4XL U3088 ( .A(\reg_file_next[8][19] ), .B(\reg_file_next[9][19] ), .C(
        \reg_file_next[10][19] ), .D(\reg_file_next[11][19] ), .S0(n2255), 
        .S1(n2243), .Y(n2508) );
  MXI4XL U3089 ( .A(\reg_file_next[8][20] ), .B(\reg_file_next[9][20] ), .C(
        \reg_file_next[10][20] ), .D(\reg_file_next[11][20] ), .S0(n2255), 
        .S1(n2250), .Y(n2516) );
  MXI4XL U3090 ( .A(\reg_file_next[8][21] ), .B(\reg_file_next[9][21] ), .C(
        \reg_file_next[10][21] ), .D(\reg_file_next[11][21] ), .S0(n2256), 
        .S1(n2248), .Y(n2524) );
  MXI4XL U3091 ( .A(\reg_file_next[8][22] ), .B(\reg_file_next[9][22] ), .C(
        \reg_file_next[10][22] ), .D(\reg_file_next[11][22] ), .S0(n2257), 
        .S1(n2251), .Y(n2532) );
  MXI4XL U3092 ( .A(\reg_file_next[8][23] ), .B(\reg_file_next[9][23] ), .C(
        \reg_file_next[10][23] ), .D(\reg_file_next[11][23] ), .S0(n2257), 
        .S1(n2244), .Y(n2540) );
  MXI4XL U3093 ( .A(\reg_file_next[8][24] ), .B(\reg_file_next[9][24] ), .C(
        \reg_file_next[10][24] ), .D(\reg_file_next[11][24] ), .S0(n2258), 
        .S1(n2244), .Y(n2548) );
  MXI4XL U3094 ( .A(\reg_file_next[8][25] ), .B(\reg_file_next[9][25] ), .C(
        \reg_file_next[10][25] ), .D(\reg_file_next[11][25] ), .S0(n2258), 
        .S1(n2245), .Y(n2556) );
  MXI4XL U3095 ( .A(\reg_file_next[8][26] ), .B(\reg_file_next[9][26] ), .C(
        \reg_file_next[10][26] ), .D(\reg_file_next[11][26] ), .S0(n2259), 
        .S1(n2245), .Y(n2564) );
  MXI4XL U3096 ( .A(\reg_file_next[8][27] ), .B(\reg_file_next[9][27] ), .C(
        \reg_file_next[10][27] ), .D(\reg_file_next[11][27] ), .S0(n2259), 
        .S1(n2245), .Y(n2572) );
  MXI4XL U3097 ( .A(\reg_file_next[8][28] ), .B(\reg_file_next[9][28] ), .C(
        \reg_file_next[10][28] ), .D(\reg_file_next[11][28] ), .S0(n2260), 
        .S1(n2246), .Y(n2580) );
  MXI4XL U3098 ( .A(\reg_file_next[8][29] ), .B(\reg_file_next[9][29] ), .C(
        \reg_file_next[10][29] ), .D(\reg_file_next[11][29] ), .S0(n2261), 
        .S1(n2246), .Y(n2588) );
  MXI4XL U3099 ( .A(\reg_file_next[8][30] ), .B(\reg_file_next[9][30] ), .C(
        \reg_file_next[10][30] ), .D(\reg_file_next[11][30] ), .S0(n2261), 
        .S1(n2246), .Y(n2596) );
  MXI4XL U3100 ( .A(\reg_file_next[8][31] ), .B(\reg_file_next[9][31] ), .C(
        \reg_file_next[10][31] ), .D(\reg_file_next[11][31] ), .S0(n2262), 
        .S1(n2250), .Y(n2604) );
  BUFX4 U3101 ( .A(n2252), .Y(n2251) );
  CLKBUFX3 U3102 ( .A(N68), .Y(n2253) );
  CLKBUFX3 U3103 ( .A(n2225), .Y(n2224) );
  CLKBUFX3 U3104 ( .A(N69), .Y(n2242) );
  CLKBUFX3 U3105 ( .A(n2247), .Y(n2252) );
  MXI2X1 U3106 ( .A(n2287), .B(n2288), .S0(N72), .Y(read_data1[0]) );
  MX4XL U3107 ( .A(n2354), .B(n2352), .C(n2353), .D(n2351), .S0(N71), .S1(N70), 
        .Y(n2288) );
  MX4XL U3108 ( .A(n2358), .B(n2356), .C(n2357), .D(n2355), .S0(N71), .S1(N70), 
        .Y(n2287) );
  MXI4XL U3109 ( .A(\reg_file_next[24][0] ), .B(\reg_file_next[25][0] ), .C(
        \reg_file_next[26][0] ), .D(\reg_file_next[27][0] ), .S0(n2267), .S1(
        n2249), .Y(n2352) );
  MXI2X1 U3110 ( .A(n2289), .B(n2290), .S0(N72), .Y(read_data1[1]) );
  MX4XL U3111 ( .A(n2362), .B(n2360), .C(n2361), .D(n2359), .S0(N71), .S1(N70), 
        .Y(n2290) );
  MX4XL U3112 ( .A(n2366), .B(n2364), .C(n2365), .D(n2363), .S0(N71), .S1(N70), 
        .Y(n2289) );
  MXI4XL U3113 ( .A(\reg_file_next[24][1] ), .B(\reg_file_next[25][1] ), .C(
        \reg_file_next[26][1] ), .D(\reg_file_next[27][1] ), .S0(n2263), .S1(
        n2248), .Y(n2360) );
  MXI2X1 U3114 ( .A(n2291), .B(n2292), .S0(N72), .Y(read_data1[2]) );
  MX4XL U3115 ( .A(n2370), .B(n2368), .C(n2369), .D(n2367), .S0(N71), .S1(N70), 
        .Y(n2292) );
  MX4XL U3116 ( .A(n2374), .B(n2372), .C(n2373), .D(n2371), .S0(N71), .S1(N70), 
        .Y(n2291) );
  MXI4XL U3117 ( .A(\reg_file_next[24][2] ), .B(\reg_file_next[25][2] ), .C(
        \reg_file_next[26][2] ), .D(\reg_file_next[27][2] ), .S0(n2263), .S1(
        n2247), .Y(n2368) );
  MXI2X1 U3118 ( .A(n2293), .B(n2294), .S0(N72), .Y(read_data1[3]) );
  MX4XL U3119 ( .A(n2378), .B(n2376), .C(n2377), .D(n2375), .S0(N71), .S1(N70), 
        .Y(n2294) );
  MX4XL U3120 ( .A(n2382), .B(n2380), .C(n2381), .D(n2379), .S0(N71), .S1(N70), 
        .Y(n2293) );
  MXI4XL U3121 ( .A(\reg_file_next[24][3] ), .B(\reg_file_next[25][3] ), .C(
        \reg_file_next[26][3] ), .D(\reg_file_next[27][3] ), .S0(n2264), .S1(
        n2247), .Y(n2376) );
  MXI2X1 U3122 ( .A(n2295), .B(n2296), .S0(N72), .Y(read_data1[4]) );
  MX4XL U3123 ( .A(n2386), .B(n2384), .C(n2385), .D(n2383), .S0(N71), .S1(N70), 
        .Y(n2296) );
  MX4XL U3124 ( .A(n2390), .B(n2388), .C(n2389), .D(n2387), .S0(N71), .S1(N70), 
        .Y(n2295) );
  MXI4XL U3125 ( .A(\reg_file_next[24][4] ), .B(\reg_file_next[25][4] ), .C(
        \reg_file_next[26][4] ), .D(\reg_file_next[27][4] ), .S0(n2264), .S1(
        n2247), .Y(n2384) );
  MXI2X1 U3126 ( .A(n2297), .B(n2298), .S0(N72), .Y(read_data1[5]) );
  MX4XL U3127 ( .A(n2394), .B(n2392), .C(n2393), .D(n2391), .S0(N71), .S1(N70), 
        .Y(n2298) );
  MX4XL U3128 ( .A(n2398), .B(n2396), .C(n2397), .D(n2395), .S0(N71), .S1(N70), 
        .Y(n2297) );
  MXI4XL U3129 ( .A(\reg_file_next[24][5] ), .B(\reg_file_next[25][5] ), .C(
        \reg_file_next[26][5] ), .D(\reg_file_next[27][5] ), .S0(n2265), .S1(
        n2248), .Y(n2392) );
  MXI2X1 U3130 ( .A(n2299), .B(n2300), .S0(N72), .Y(read_data1[6]) );
  MX4XL U3131 ( .A(n2402), .B(n2400), .C(n2401), .D(n2399), .S0(N71), .S1(N70), 
        .Y(n2300) );
  MX4XL U3132 ( .A(n2406), .B(n2404), .C(n2405), .D(n2403), .S0(N71), .S1(N70), 
        .Y(n2299) );
  MXI4XL U3133 ( .A(\reg_file_next[24][6] ), .B(\reg_file_next[25][6] ), .C(
        \reg_file_next[26][6] ), .D(\reg_file_next[27][6] ), .S0(n2265), .S1(
        n2248), .Y(n2400) );
  MXI2X1 U3134 ( .A(n2301), .B(n2302), .S0(N72), .Y(read_data1[7]) );
  MX4XL U3135 ( .A(n2410), .B(n2408), .C(n2409), .D(n2407), .S0(N71), .S1(N70), 
        .Y(n2302) );
  MX4XL U3136 ( .A(n2414), .B(n2412), .C(n2413), .D(n2411), .S0(N71), .S1(N70), 
        .Y(n2301) );
  MXI4XL U3137 ( .A(\reg_file_next[24][7] ), .B(\reg_file_next[25][7] ), .C(
        \reg_file_next[26][7] ), .D(\reg_file_next[27][7] ), .S0(n2266), .S1(
        n2249), .Y(n2408) );
  MXI2X1 U3138 ( .A(n2303), .B(n2304), .S0(N72), .Y(read_data1[8]) );
  MX4XL U3139 ( .A(n2418), .B(n2416), .C(n2417), .D(n2415), .S0(N71), .S1(N70), 
        .Y(n2304) );
  MX4XL U3140 ( .A(n2422), .B(n2420), .C(n2421), .D(n2419), .S0(N71), .S1(N70), 
        .Y(n2303) );
  MXI4XL U3141 ( .A(\reg_file_next[24][8] ), .B(\reg_file_next[25][8] ), .C(
        \reg_file_next[26][8] ), .D(\reg_file_next[27][8] ), .S0(n2267), .S1(
        n2249), .Y(n2416) );
  MXI2X1 U3142 ( .A(n2305), .B(n2306), .S0(N72), .Y(read_data1[9]) );
  MX4XL U3143 ( .A(n2426), .B(n2424), .C(n2425), .D(n2423), .S0(N71), .S1(N70), 
        .Y(n2306) );
  MX4XL U3144 ( .A(n2430), .B(n2428), .C(n2429), .D(n2427), .S0(N71), .S1(N70), 
        .Y(n2305) );
  MXI4XL U3145 ( .A(\reg_file_next[24][9] ), .B(\reg_file_next[25][9] ), .C(
        \reg_file_next[26][9] ), .D(\reg_file_next[27][9] ), .S0(n2267), .S1(
        n2249), .Y(n2424) );
  MXI2X1 U3146 ( .A(n2307), .B(n2308), .S0(N72), .Y(read_data1[10]) );
  MX4XL U3147 ( .A(n2434), .B(n2432), .C(n2433), .D(n2431), .S0(N71), .S1(N70), 
        .Y(n2308) );
  MX4XL U3148 ( .A(n2438), .B(n2436), .C(n2437), .D(n2435), .S0(N71), .S1(N70), 
        .Y(n2307) );
  MXI4XL U3149 ( .A(\reg_file_next[24][10] ), .B(\reg_file_next[25][10] ), .C(
        \reg_file_next[26][10] ), .D(\reg_file_next[27][10] ), .S0(n2268), 
        .S1(n2250), .Y(n2432) );
  MXI2X1 U3150 ( .A(n2309), .B(n2310), .S0(N72), .Y(read_data1[11]) );
  MX4XL U3151 ( .A(n2442), .B(n2440), .C(n2441), .D(n2439), .S0(N71), .S1(N70), 
        .Y(n2310) );
  MX4XL U3152 ( .A(n2446), .B(n2444), .C(n2445), .D(n2443), .S0(N71), .S1(N70), 
        .Y(n2309) );
  MXI4XL U3153 ( .A(\reg_file_next[24][11] ), .B(\reg_file_next[25][11] ), .C(
        \reg_file_next[26][11] ), .D(\reg_file_next[27][11] ), .S0(n2268), 
        .S1(n2250), .Y(n2440) );
  MXI2X1 U3154 ( .A(n2311), .B(n2312), .S0(N72), .Y(read_data1[12]) );
  MX4XL U3155 ( .A(n2450), .B(n2448), .C(n2449), .D(n2447), .S0(N71), .S1(N70), 
        .Y(n2312) );
  MX4XL U3156 ( .A(n2454), .B(n2452), .C(n2453), .D(n2451), .S0(N71), .S1(N70), 
        .Y(n2311) );
  MXI4XL U3157 ( .A(\reg_file_next[24][12] ), .B(\reg_file_next[25][12] ), .C(
        \reg_file_next[26][12] ), .D(\reg_file_next[27][12] ), .S0(n2269), 
        .S1(n2251), .Y(n2448) );
  MXI2X1 U3158 ( .A(n2313), .B(n2314), .S0(N72), .Y(read_data1[13]) );
  MX4XL U3159 ( .A(n2458), .B(n2456), .C(n2457), .D(n2455), .S0(N71), .S1(N70), 
        .Y(n2314) );
  MX4XL U3160 ( .A(n2462), .B(n2460), .C(n2461), .D(n2459), .S0(N71), .S1(N70), 
        .Y(n2313) );
  MXI4XL U3161 ( .A(\reg_file_next[24][13] ), .B(\reg_file_next[25][13] ), .C(
        \reg_file_next[26][13] ), .D(\reg_file_next[27][13] ), .S0(n2269), 
        .S1(n2251), .Y(n2456) );
  MXI2X1 U3162 ( .A(n2315), .B(n2316), .S0(N72), .Y(read_data1[14]) );
  MX4XL U3163 ( .A(n2466), .B(n2464), .C(n2465), .D(n2463), .S0(N71), .S1(N70), 
        .Y(n2316) );
  MX4XL U3164 ( .A(n2470), .B(n2468), .C(n2469), .D(n2467), .S0(N71), .S1(N70), 
        .Y(n2315) );
  MXI4XL U3165 ( .A(\reg_file_next[24][14] ), .B(\reg_file_next[25][14] ), .C(
        \reg_file_next[26][14] ), .D(\reg_file_next[27][14] ), .S0(n2270), 
        .S1(n2251), .Y(n2464) );
  MXI2X1 U3166 ( .A(n2317), .B(n2318), .S0(N72), .Y(read_data1[15]) );
  MX4XL U3167 ( .A(n2474), .B(n2472), .C(n2473), .D(n2471), .S0(N71), .S1(N70), 
        .Y(n2318) );
  MX4XL U3168 ( .A(n2478), .B(n2476), .C(n2477), .D(n2475), .S0(N71), .S1(N70), 
        .Y(n2317) );
  MXI4XL U3169 ( .A(\reg_file_next[24][15] ), .B(\reg_file_next[25][15] ), .C(
        \reg_file_next[26][15] ), .D(\reg_file_next[27][15] ), .S0(n2267), 
        .S1(n2252), .Y(n2472) );
  MXI2X1 U3170 ( .A(n2319), .B(n2320), .S0(N72), .Y(read_data1[16]) );
  MX4XL U3171 ( .A(n2482), .B(n2480), .C(n2481), .D(n2479), .S0(N71), .S1(N70), 
        .Y(n2320) );
  MX4XL U3172 ( .A(n2486), .B(n2484), .C(n2485), .D(n2483), .S0(N71), .S1(N70), 
        .Y(n2319) );
  MXI4XL U3173 ( .A(\reg_file_next[24][16] ), .B(\reg_file_next[25][16] ), .C(
        \reg_file_next[26][16] ), .D(\reg_file_next[27][16] ), .S0(n2253), 
        .S1(n2242), .Y(n2480) );
  MXI2X1 U3174 ( .A(n2321), .B(n2322), .S0(N72), .Y(read_data1[17]) );
  MX4XL U3175 ( .A(n2490), .B(n2488), .C(n2489), .D(n2487), .S0(N71), .S1(N70), 
        .Y(n2322) );
  MX4XL U3176 ( .A(n2494), .B(n2492), .C(n2493), .D(n2491), .S0(N71), .S1(N70), 
        .Y(n2321) );
  MXI4XL U3177 ( .A(\reg_file_next[24][17] ), .B(\reg_file_next[25][17] ), .C(
        \reg_file_next[26][17] ), .D(\reg_file_next[27][17] ), .S0(n2253), 
        .S1(n2242), .Y(n2488) );
  MXI2X1 U3178 ( .A(n2323), .B(n2324), .S0(N72), .Y(read_data1[18]) );
  MX4XL U3179 ( .A(n2498), .B(n2496), .C(n2497), .D(n2495), .S0(N71), .S1(N70), 
        .Y(n2324) );
  MX4XL U3180 ( .A(n2502), .B(n2500), .C(n2501), .D(n2499), .S0(N71), .S1(N70), 
        .Y(n2323) );
  MXI4XL U3181 ( .A(\reg_file_next[24][18] ), .B(\reg_file_next[25][18] ), .C(
        \reg_file_next[26][18] ), .D(\reg_file_next[27][18] ), .S0(n2254), 
        .S1(n2243), .Y(n2496) );
  MXI2X1 U3182 ( .A(n2325), .B(n2326), .S0(N72), .Y(read_data1[19]) );
  MX4XL U3183 ( .A(n2506), .B(n2504), .C(n2505), .D(n2503), .S0(N71), .S1(N70), 
        .Y(n2326) );
  MX4XL U3184 ( .A(n2510), .B(n2508), .C(n2509), .D(n2507), .S0(N71), .S1(N70), 
        .Y(n2325) );
  MXI4XL U3185 ( .A(\reg_file_next[24][19] ), .B(\reg_file_next[25][19] ), .C(
        \reg_file_next[26][19] ), .D(\reg_file_next[27][19] ), .S0(n2255), 
        .S1(n2243), .Y(n2504) );
  MXI2X1 U3186 ( .A(n2327), .B(n2328), .S0(N72), .Y(read_data1[20]) );
  MX4XL U3187 ( .A(n2514), .B(n2512), .C(n2513), .D(n2511), .S0(N71), .S1(N70), 
        .Y(n2328) );
  MX4XL U3188 ( .A(n2518), .B(n2516), .C(n2517), .D(n2515), .S0(N71), .S1(N70), 
        .Y(n2327) );
  MXI4XL U3189 ( .A(\reg_file_next[24][20] ), .B(\reg_file_next[25][20] ), .C(
        \reg_file_next[26][20] ), .D(\reg_file_next[27][20] ), .S0(n2255), 
        .S1(n2243), .Y(n2512) );
  MXI2X1 U3190 ( .A(n2329), .B(n2330), .S0(N72), .Y(read_data1[21]) );
  MX4XL U3191 ( .A(n2522), .B(n2520), .C(n2521), .D(n2519), .S0(N71), .S1(N70), 
        .Y(n2330) );
  MX4XL U3192 ( .A(n2526), .B(n2524), .C(n2525), .D(n2523), .S0(N71), .S1(N70), 
        .Y(n2329) );
  MXI4XL U3193 ( .A(\reg_file_next[24][21] ), .B(\reg_file_next[25][21] ), .C(
        \reg_file_next[26][21] ), .D(\reg_file_next[27][21] ), .S0(n2256), 
        .S1(n2243), .Y(n2520) );
  MXI2X1 U3194 ( .A(n2331), .B(n2332), .S0(N72), .Y(read_data1[22]) );
  MX4XL U3195 ( .A(n2530), .B(n2528), .C(n2529), .D(n2527), .S0(N71), .S1(N70), 
        .Y(n2332) );
  MX4XL U3196 ( .A(n2534), .B(n2532), .C(n2533), .D(n2531), .S0(N71), .S1(N70), 
        .Y(n2331) );
  MXI4XL U3197 ( .A(\reg_file_next[24][22] ), .B(\reg_file_next[25][22] ), .C(
        \reg_file_next[26][22] ), .D(\reg_file_next[27][22] ), .S0(n2256), 
        .S1(n2247), .Y(n2528) );
  MXI2X1 U3198 ( .A(n2333), .B(n2334), .S0(N72), .Y(read_data1[23]) );
  MX4XL U3199 ( .A(n2538), .B(n2536), .C(n2537), .D(n2535), .S0(N71), .S1(N70), 
        .Y(n2334) );
  MX4XL U3200 ( .A(n2542), .B(n2540), .C(n2541), .D(n2539), .S0(N71), .S1(N70), 
        .Y(n2333) );
  MXI4XL U3201 ( .A(\reg_file_next[24][23] ), .B(\reg_file_next[25][23] ), .C(
        \reg_file_next[26][23] ), .D(\reg_file_next[27][23] ), .S0(n2257), 
        .S1(n2244), .Y(n2536) );
  MXI2X1 U3202 ( .A(n2335), .B(n2336), .S0(N72), .Y(read_data1[24]) );
  MX4XL U3203 ( .A(n2546), .B(n2544), .C(n2545), .D(n2543), .S0(N71), .S1(N70), 
        .Y(n2336) );
  MX4XL U3204 ( .A(n2550), .B(n2548), .C(n2549), .D(n2547), .S0(N71), .S1(N70), 
        .Y(n2335) );
  MXI4XL U3205 ( .A(\reg_file_next[24][24] ), .B(\reg_file_next[25][24] ), .C(
        \reg_file_next[26][24] ), .D(\reg_file_next[27][24] ), .S0(n2257), 
        .S1(n2244), .Y(n2544) );
  MXI2X1 U3206 ( .A(n2337), .B(n2338), .S0(N72), .Y(read_data1[25]) );
  MX4XL U3207 ( .A(n2554), .B(n2552), .C(n2553), .D(n2551), .S0(N71), .S1(N70), 
        .Y(n2338) );
  MX4XL U3208 ( .A(n2558), .B(n2556), .C(n2557), .D(n2555), .S0(N71), .S1(N70), 
        .Y(n2337) );
  MXI4XL U3209 ( .A(\reg_file_next[24][25] ), .B(\reg_file_next[25][25] ), .C(
        \reg_file_next[26][25] ), .D(\reg_file_next[27][25] ), .S0(n2258), 
        .S1(n2244), .Y(n2552) );
  MXI2X1 U3210 ( .A(n2339), .B(n2340), .S0(N72), .Y(read_data1[26]) );
  MX4XL U3211 ( .A(n2562), .B(n2560), .C(n2561), .D(n2559), .S0(N71), .S1(N70), 
        .Y(n2340) );
  MX4XL U3212 ( .A(n2566), .B(n2564), .C(n2565), .D(n2563), .S0(N71), .S1(N70), 
        .Y(n2339) );
  MXI4XL U3213 ( .A(\reg_file_next[24][26] ), .B(\reg_file_next[25][26] ), .C(
        \reg_file_next[26][26] ), .D(\reg_file_next[27][26] ), .S0(n2259), 
        .S1(n2245), .Y(n2560) );
  MXI2X1 U3214 ( .A(n2341), .B(n2342), .S0(N72), .Y(read_data1[27]) );
  MX4XL U3215 ( .A(n2570), .B(n2568), .C(n2569), .D(n2567), .S0(N71), .S1(N70), 
        .Y(n2342) );
  MX4XL U3216 ( .A(n2574), .B(n2572), .C(n2573), .D(n2571), .S0(N71), .S1(N70), 
        .Y(n2341) );
  MXI4XL U3217 ( .A(\reg_file_next[24][27] ), .B(\reg_file_next[25][27] ), .C(
        \reg_file_next[26][27] ), .D(\reg_file_next[27][27] ), .S0(n2259), 
        .S1(n2245), .Y(n2568) );
  MXI2X1 U3218 ( .A(n2343), .B(n2344), .S0(N72), .Y(read_data1[28]) );
  MX4XL U3219 ( .A(n2578), .B(n2576), .C(n2577), .D(n2575), .S0(N71), .S1(N70), 
        .Y(n2344) );
  MX4XL U3220 ( .A(n2582), .B(n2580), .C(n2581), .D(n2579), .S0(N71), .S1(N70), 
        .Y(n2343) );
  MXI4XL U3221 ( .A(\reg_file_next[24][28] ), .B(\reg_file_next[25][28] ), .C(
        \reg_file_next[26][28] ), .D(\reg_file_next[27][28] ), .S0(n2260), 
        .S1(n2245), .Y(n2576) );
  MXI2X1 U3222 ( .A(n2345), .B(n2346), .S0(N72), .Y(read_data1[29]) );
  MX4XL U3223 ( .A(n2586), .B(n2584), .C(n2585), .D(n2583), .S0(N71), .S1(N70), 
        .Y(n2346) );
  MX4XL U3224 ( .A(n2590), .B(n2588), .C(n2589), .D(n2587), .S0(N71), .S1(N70), 
        .Y(n2345) );
  MXI4XL U3225 ( .A(\reg_file_next[24][29] ), .B(\reg_file_next[25][29] ), .C(
        \reg_file_next[26][29] ), .D(\reg_file_next[27][29] ), .S0(n2260), 
        .S1(n2246), .Y(n2584) );
  MXI2X1 U3226 ( .A(n2347), .B(n2348), .S0(N72), .Y(read_data1[30]) );
  MX4XL U3227 ( .A(n2594), .B(n2592), .C(n2593), .D(n2591), .S0(N71), .S1(N70), 
        .Y(n2348) );
  MX4XL U3228 ( .A(n2598), .B(n2596), .C(n2597), .D(n2595), .S0(N71), .S1(N70), 
        .Y(n2347) );
  MXI4XL U3229 ( .A(\reg_file_next[24][30] ), .B(\reg_file_next[25][30] ), .C(
        \reg_file_next[26][30] ), .D(\reg_file_next[27][30] ), .S0(n2261), 
        .S1(n2246), .Y(n2592) );
  MXI2X1 U3230 ( .A(n2349), .B(n2350), .S0(N72), .Y(read_data1[31]) );
  MX4XL U3231 ( .A(n2602), .B(n2600), .C(n2601), .D(n2599), .S0(N71), .S1(N70), 
        .Y(n2350) );
  MX4XL U3232 ( .A(n2606), .B(n2604), .C(n2605), .D(n2603), .S0(N71), .S1(N70), 
        .Y(n2349) );
  MXI4XL U3233 ( .A(\reg_file_next[24][31] ), .B(\reg_file_next[25][31] ), .C(
        \reg_file_next[26][31] ), .D(\reg_file_next[27][31] ), .S0(n2261), 
        .S1(n2251), .Y(n2600) );
  MXI2XL U3234 ( .A(n2607), .B(n2608), .S0(N77), .Y(read_data2[0]) );
  MX4XL U3235 ( .A(n2674), .B(n2672), .C(n2673), .D(n2671), .S0(N76), .S1(N75), 
        .Y(n2608) );
  MX4XL U3236 ( .A(n2678), .B(n2676), .C(n2677), .D(n2675), .S0(N76), .S1(N75), 
        .Y(n2607) );
  MXI4XL U3237 ( .A(\reg_file_next[24][0] ), .B(\reg_file_next[25][0] ), .C(
        \reg_file_next[26][0] ), .D(\reg_file_next[27][0] ), .S0(n2238), .S1(
        n2219), .Y(n2672) );
  MXI2XL U3238 ( .A(n2609), .B(n2610), .S0(N77), .Y(read_data2[1]) );
  MX4XL U3239 ( .A(n2682), .B(n2680), .C(n2681), .D(n2679), .S0(N76), .S1(N75), 
        .Y(n2610) );
  MX4XL U3240 ( .A(n2686), .B(n2684), .C(n2685), .D(n2683), .S0(N76), .S1(N75), 
        .Y(n2609) );
  MXI4XL U3241 ( .A(\reg_file_next[24][1] ), .B(\reg_file_next[25][1] ), .C(
        \reg_file_next[26][1] ), .D(\reg_file_next[27][1] ), .S0(n2234), .S1(
        n2217), .Y(n2680) );
  MXI2XL U3242 ( .A(n2611), .B(n2612), .S0(N77), .Y(read_data2[2]) );
  MX4XL U3243 ( .A(n2690), .B(n2688), .C(n2689), .D(n2687), .S0(N76), .S1(N75), 
        .Y(n2612) );
  MX4XL U3244 ( .A(n2694), .B(n2692), .C(n2693), .D(n2691), .S0(N76), .S1(N75), 
        .Y(n2611) );
  MXI4XL U3245 ( .A(\reg_file_next[24][2] ), .B(\reg_file_next[25][2] ), .C(
        \reg_file_next[26][2] ), .D(\reg_file_next[27][2] ), .S0(n2234), .S1(
        n2217), .Y(n2688) );
  MXI2XL U3246 ( .A(n2613), .B(n2614), .S0(N77), .Y(read_data2[3]) );
  MX4XL U3247 ( .A(n2698), .B(n2696), .C(n2697), .D(n2695), .S0(N76), .S1(N75), 
        .Y(n2614) );
  MX4XL U3248 ( .A(n2702), .B(n2700), .C(n2701), .D(n2699), .S0(N76), .S1(N75), 
        .Y(n2613) );
  MXI4XL U3249 ( .A(\reg_file_next[24][3] ), .B(\reg_file_next[25][3] ), .C(
        \reg_file_next[26][3] ), .D(\reg_file_next[27][3] ), .S0(n2235), .S1(
        n2217), .Y(n2696) );
  MXI2XL U3250 ( .A(n2615), .B(n2616), .S0(N77), .Y(read_data2[4]) );
  MX4XL U3251 ( .A(n2706), .B(n2704), .C(n2705), .D(n2703), .S0(N76), .S1(N75), 
        .Y(n2616) );
  MX4XL U3252 ( .A(n2710), .B(n2708), .C(n2709), .D(n2707), .S0(N76), .S1(N75), 
        .Y(n2615) );
  MXI4XL U3253 ( .A(\reg_file_next[24][4] ), .B(\reg_file_next[25][4] ), .C(
        \reg_file_next[26][4] ), .D(\reg_file_next[27][4] ), .S0(n2235), .S1(
        n2218), .Y(n2704) );
  MXI2XL U3254 ( .A(n2617), .B(n2618), .S0(N77), .Y(read_data2[5]) );
  MX4XL U3255 ( .A(n2714), .B(n2712), .C(n2713), .D(n2711), .S0(N76), .S1(N75), 
        .Y(n2618) );
  MX4XL U3256 ( .A(n2718), .B(n2716), .C(n2717), .D(n2715), .S0(N76), .S1(N75), 
        .Y(n2617) );
  MXI4XL U3257 ( .A(\reg_file_next[24][5] ), .B(\reg_file_next[25][5] ), .C(
        \reg_file_next[26][5] ), .D(\reg_file_next[27][5] ), .S0(n2236), .S1(
        n2218), .Y(n2712) );
  MX4XL U3258 ( .A(n2722), .B(n2720), .C(n2721), .D(n2719), .S0(N76), .S1(N75), 
        .Y(n2620) );
  MX4XL U3259 ( .A(n2726), .B(n2724), .C(n2725), .D(n2723), .S0(N76), .S1(N75), 
        .Y(n2619) );
  MX4XL U3260 ( .A(n2730), .B(n2728), .C(n2729), .D(n2727), .S0(N76), .S1(N75), 
        .Y(n2622) );
  MX4XL U3261 ( .A(n2734), .B(n2732), .C(n2733), .D(n2731), .S0(N76), .S1(N75), 
        .Y(n2621) );
  MX4XL U3262 ( .A(n2738), .B(n2736), .C(n2737), .D(n2735), .S0(N76), .S1(N75), 
        .Y(n2624) );
  MX4XL U3263 ( .A(n2742), .B(n2740), .C(n2741), .D(n2739), .S0(N76), .S1(N75), 
        .Y(n2623) );
  MX4XL U3264 ( .A(n2746), .B(n2744), .C(n2745), .D(n2743), .S0(N76), .S1(N75), 
        .Y(n2626) );
  MX4XL U3265 ( .A(n2750), .B(n2748), .C(n2749), .D(n2747), .S0(N76), .S1(N75), 
        .Y(n2625) );
  MX4XL U3266 ( .A(n2754), .B(n2752), .C(n2753), .D(n2751), .S0(N76), .S1(N75), 
        .Y(n2628) );
  MX4XL U3267 ( .A(n2758), .B(n2756), .C(n2757), .D(n2755), .S0(N76), .S1(N75), 
        .Y(n2627) );
  MX4XL U3268 ( .A(n2762), .B(n2760), .C(n2761), .D(n2759), .S0(N76), .S1(N75), 
        .Y(n2630) );
  MX4XL U3269 ( .A(n2766), .B(n2764), .C(n2765), .D(n2763), .S0(N76), .S1(N75), 
        .Y(n2629) );
  MX4XL U3270 ( .A(n2770), .B(n2768), .C(n2769), .D(n2767), .S0(N76), .S1(N75), 
        .Y(n2632) );
  MX4XL U3271 ( .A(n2774), .B(n2772), .C(n2773), .D(n2771), .S0(N76), .S1(N75), 
        .Y(n2631) );
  MX4XL U3272 ( .A(n2778), .B(n2776), .C(n2777), .D(n2775), .S0(N76), .S1(N75), 
        .Y(n2634) );
  MX4XL U3273 ( .A(n2782), .B(n2780), .C(n2781), .D(n2779), .S0(N76), .S1(N75), 
        .Y(n2633) );
  MX4XL U3274 ( .A(n2786), .B(n2784), .C(n2785), .D(n2783), .S0(N76), .S1(N75), 
        .Y(n2636) );
  MX4XL U3275 ( .A(n2790), .B(n2788), .C(n2789), .D(n2787), .S0(N76), .S1(N75), 
        .Y(n2635) );
  MX4XL U3276 ( .A(n2794), .B(n2792), .C(n2793), .D(n2791), .S0(N76), .S1(N75), 
        .Y(n2638) );
  MX4XL U3277 ( .A(n2798), .B(n2796), .C(n2797), .D(n2795), .S0(N76), .S1(N75), 
        .Y(n2637) );
  MX4XL U3278 ( .A(n2802), .B(n2800), .C(n2801), .D(n2799), .S0(N76), .S1(N75), 
        .Y(n2640) );
  MX4XL U3279 ( .A(n2806), .B(n2804), .C(n2805), .D(n2803), .S0(N76), .S1(N75), 
        .Y(n2639) );
  MX4XL U3280 ( .A(n2810), .B(n2808), .C(n2809), .D(n2807), .S0(N76), .S1(N75), 
        .Y(n2642) );
  MX4XL U3281 ( .A(n2814), .B(n2812), .C(n2813), .D(n2811), .S0(N76), .S1(N75), 
        .Y(n2641) );
  MX4XL U3282 ( .A(n2818), .B(n2816), .C(n2817), .D(n2815), .S0(N76), .S1(N75), 
        .Y(n2644) );
  MX4XL U3283 ( .A(n2822), .B(n2820), .C(n2821), .D(n2819), .S0(N76), .S1(N75), 
        .Y(n2643) );
  MX4XL U3284 ( .A(n2826), .B(n2824), .C(n2825), .D(n2823), .S0(N76), .S1(N75), 
        .Y(n2646) );
  MX4XL U3285 ( .A(n2830), .B(n2828), .C(n2829), .D(n2827), .S0(N76), .S1(N75), 
        .Y(n2645) );
  MX4XL U3286 ( .A(n2834), .B(n2832), .C(n2833), .D(n2831), .S0(N76), .S1(N75), 
        .Y(n2648) );
  MX4XL U3287 ( .A(n2838), .B(n2836), .C(n2837), .D(n2835), .S0(N76), .S1(N75), 
        .Y(n2647) );
  MX4XL U3288 ( .A(n2842), .B(n2840), .C(n2841), .D(n2839), .S0(N76), .S1(N75), 
        .Y(n2650) );
  MX4XL U3289 ( .A(n2846), .B(n2844), .C(n2845), .D(n2843), .S0(N76), .S1(N75), 
        .Y(n2649) );
  MX4XL U3290 ( .A(n2850), .B(n2848), .C(n2849), .D(n2847), .S0(N76), .S1(N75), 
        .Y(n2652) );
  MX4XL U3291 ( .A(n2854), .B(n2852), .C(n2853), .D(n2851), .S0(N76), .S1(N75), 
        .Y(n2651) );
  MX4XL U3292 ( .A(n2858), .B(n2856), .C(n2857), .D(n2855), .S0(N76), .S1(N75), 
        .Y(n2654) );
  MX4XL U3293 ( .A(n2862), .B(n2860), .C(n2861), .D(n2859), .S0(N76), .S1(N75), 
        .Y(n2653) );
  MX4XL U3294 ( .A(n2866), .B(n2864), .C(n2865), .D(n2863), .S0(N76), .S1(N75), 
        .Y(n2656) );
  MX4XL U3295 ( .A(n2870), .B(n2868), .C(n2869), .D(n2867), .S0(N76), .S1(N75), 
        .Y(n2655) );
  MX4XL U3296 ( .A(n2874), .B(n2872), .C(n2873), .D(n2871), .S0(N76), .S1(N75), 
        .Y(n2658) );
  MX4XL U3297 ( .A(n2878), .B(n2876), .C(n2877), .D(n2875), .S0(N76), .S1(N75), 
        .Y(n2657) );
  MX4XL U3298 ( .A(n2882), .B(n2880), .C(n2881), .D(n2879), .S0(N76), .S1(N75), 
        .Y(n2660) );
  MX4XL U3299 ( .A(n2886), .B(n2884), .C(n2885), .D(n2883), .S0(N76), .S1(N75), 
        .Y(n2659) );
  MX4XL U3300 ( .A(n2890), .B(n2888), .C(n2889), .D(n2887), .S0(N76), .S1(N75), 
        .Y(n2662) );
  MX4XL U3301 ( .A(n2894), .B(n2892), .C(n2893), .D(n2891), .S0(N76), .S1(N75), 
        .Y(n2661) );
  MX4XL U3302 ( .A(n2898), .B(n2896), .C(n2897), .D(n2895), .S0(N76), .S1(N75), 
        .Y(n2664) );
  MX4XL U3303 ( .A(n2902), .B(n2900), .C(n2901), .D(n2899), .S0(N76), .S1(N75), 
        .Y(n2663) );
  MX4XL U3304 ( .A(n2906), .B(n2904), .C(n2905), .D(n2903), .S0(N76), .S1(N75), 
        .Y(n2666) );
  MX4XL U3305 ( .A(n2910), .B(n2908), .C(n2909), .D(n2907), .S0(N76), .S1(N75), 
        .Y(n2665) );
  MX4XL U3306 ( .A(n2914), .B(n2912), .C(n2913), .D(n2911), .S0(N76), .S1(N75), 
        .Y(n2668) );
  MX4XL U3307 ( .A(n2918), .B(n2916), .C(n2917), .D(n2915), .S0(N76), .S1(N75), 
        .Y(n2667) );
  MX4XL U3308 ( .A(n2922), .B(n2920), .C(n2921), .D(n2919), .S0(N76), .S1(N75), 
        .Y(n2670) );
  MX4XL U3309 ( .A(n2926), .B(n2924), .C(n2925), .D(n2923), .S0(N76), .S1(N75), 
        .Y(n2669) );
  CLKBUFX3 U3310 ( .A(N74), .Y(n2223) );
  CLKBUFX3 U3311 ( .A(rst_n), .Y(n2286) );
  CLKINVX1 U3312 ( .A(ICACHE_stall), .Y(n70) );
  CLKINVX1 U3313 ( .A(n3025), .Y(n31) );
  AOI221XL U3314 ( .A0(EX_Rt[4]), .A1(n3026), .B0(EX_Rd[4]), .B1(n3027), .C0(
        n3028), .Y(n3025) );
  CLKINVX1 U3315 ( .A(n3029), .Y(n30) );
  AOI221XL U3316 ( .A0(EX_Rt[3]), .A1(n3026), .B0(EX_Rd[3]), .B1(n3027), .C0(
        n3028), .Y(n3029) );
  CLKINVX1 U3317 ( .A(n3030), .Y(n29) );
  AOI221XL U3318 ( .A0(EX_Rt[2]), .A1(n3026), .B0(EX_Rd[2]), .B1(n3027), .C0(
        n3028), .Y(n3030) );
  CLKINVX1 U3319 ( .A(n3031), .Y(n28) );
  AOI221XL U3320 ( .A0(EX_Rt[1]), .A1(n3026), .B0(EX_Rd[1]), .B1(n3027), .C0(
        n3028), .Y(n3031) );
  CLKINVX1 U3321 ( .A(n3032), .Y(n27) );
  AOI221XL U3322 ( .A0(EX_Rt[0]), .A1(n3026), .B0(EX_Rd[0]), .B1(n3027), .C0(
        n3028), .Y(n3032) );
  AND2X1 U3323 ( .A(EX_reg[5]), .B(n3026), .Y(n3028) );
  NOR2X1 U3324 ( .A(n3026), .B(EX_reg[5]), .Y(n3027) );
  OAI211X1 U3325 ( .A0(n3249), .A1(n2139), .B0(n3039), .C0(n3040), .Y(n1352)
         );
  AOI222XL U3326 ( .A0(read_data1[2]), .A1(n2132), .B0(PC_plus4[2]), .B1(n3035), .C0(InstReg[0]), .C1(n2131), .Y(n3040) );
  NAND2X1 U3327 ( .A(BranchAddr[2]), .B(n3036), .Y(n3039) );
  AOI222XL U3328 ( .A0(read_data1[3]), .A1(n2132), .B0(PC_plus4[3]), .B1(n3035), .C0(InstReg[1]), .C1(n2131), .Y(n3042) );
  AOI222XL U3329 ( .A0(read_data1[4]), .A1(n2132), .B0(PC_plus4[4]), .B1(n3035), .C0(InstReg[2]), .C1(n2131), .Y(n3044) );
  AOI222XL U3330 ( .A0(read_data1[5]), .A1(n2132), .B0(PC_plus4[5]), .B1(n3035), .C0(InstReg[3]), .C1(n2131), .Y(n3046) );
  AOI222XL U3331 ( .A0(read_data1[6]), .A1(n2132), .B0(PC_plus4[6]), .B1(n3035), .C0(InstReg[4]), .C1(n2131), .Y(n3048) );
  AOI222XL U3332 ( .A0(read_data1[7]), .A1(n2132), .B0(PC_plus4[7]), .B1(n3035), .C0(InstReg[5]), .C1(n2131), .Y(n3050) );
  AOI222XL U3333 ( .A0(read_data1[8]), .A1(n2132), .B0(PC_plus4[8]), .B1(n3035), .C0(InstReg[6]), .C1(n2131), .Y(n3052) );
  AOI222XL U3334 ( .A0(read_data1[9]), .A1(n2132), .B0(PC_plus4[9]), .B1(n3035), .C0(InstReg[7]), .C1(n2131), .Y(n3054) );
  AOI222XL U3335 ( .A0(read_data1[10]), .A1(n2132), .B0(PC_plus4[10]), .B1(
        n3035), .C0(InstReg[8]), .C1(n2131), .Y(n3056) );
  AOI222XL U3336 ( .A0(read_data1[11]), .A1(n2132), .B0(PC_plus4[11]), .B1(
        n3035), .C0(InstReg[9]), .C1(n2131), .Y(n3058) );
  AOI222XL U3337 ( .A0(read_data1[12]), .A1(n2132), .B0(PC_plus4[12]), .B1(
        n3035), .C0(InstReg[10]), .C1(n2131), .Y(n3060) );
  AOI222XL U3338 ( .A0(read_data1[13]), .A1(n2132), .B0(PC_plus4[13]), .B1(
        n3035), .C0(InstReg[11]), .C1(n2131), .Y(n3062) );
  AOI222XL U3339 ( .A0(read_data1[14]), .A1(n2132), .B0(PC_plus4[14]), .B1(
        n3035), .C0(InstReg[12]), .C1(n2131), .Y(n3064) );
  AOI222XL U3340 ( .A0(read_data1[15]), .A1(n2132), .B0(PC_plus4[15]), .B1(
        n3035), .C0(InstReg[13]), .C1(n2131), .Y(n3066) );
  AOI222XL U3341 ( .A0(read_data1[16]), .A1(n2132), .B0(PC_plus4[16]), .B1(
        n3035), .C0(InstReg[14]), .C1(n2131), .Y(n3068) );
  AOI222XL U3342 ( .A0(read_data1[17]), .A1(n2132), .B0(PC_plus4[17]), .B1(
        n3035), .C0(InstReg[15]), .C1(n2131), .Y(n3070) );
  AOI222XL U3343 ( .A0(read_data1[18]), .A1(n2132), .B0(PC_plus4[18]), .B1(
        n3035), .C0(n2226), .C1(n2131), .Y(n3072) );
  AOI222XL U3344 ( .A0(read_data1[19]), .A1(n2132), .B0(PC_plus4[19]), .B1(
        n3035), .C0(n2223), .C1(n2131), .Y(n3074) );
  AOI222XL U3345 ( .A0(read_data1[20]), .A1(n2132), .B0(PC_plus4[20]), .B1(
        n3035), .C0(N75), .C1(n2131), .Y(n3076) );
  AOI222XL U3346 ( .A0(read_data1[21]), .A1(n2132), .B0(PC_plus4[21]), .B1(
        n3035), .C0(N76), .C1(n2131), .Y(n3078) );
  AOI222XL U3347 ( .A0(read_data1[22]), .A1(n2132), .B0(PC_plus4[22]), .B1(
        n3035), .C0(N77), .C1(n2131), .Y(n3080) );
  AOI222XL U3348 ( .A0(read_data1[23]), .A1(n2132), .B0(PC_plus4[23]), .B1(
        n3035), .C0(n2264), .C1(n2131), .Y(n3082) );
  AOI222XL U3349 ( .A0(read_data1[24]), .A1(n2132), .B0(PC_plus4[24]), .B1(
        n3035), .C0(n2252), .C1(n2131), .Y(n3084) );
  AOI222XL U3350 ( .A0(read_data1[25]), .A1(n2132), .B0(PC_plus4[25]), .B1(
        n3035), .C0(N70), .C1(n2131), .Y(n3086) );
  AOI222XL U3351 ( .A0(read_data1[26]), .A1(n2132), .B0(PC_plus4[26]), .B1(
        n3035), .C0(N71), .C1(n2131), .Y(n3088) );
  AOI222XL U3352 ( .A0(read_data1[27]), .A1(n2132), .B0(PC_plus4[27]), .B1(
        n3035), .C0(N72), .C1(n2131), .Y(n3090) );
  AOI222XL U3353 ( .A0(read_data1[28]), .A1(n2132), .B0(PC_plus4[28]), .B1(
        n3035), .C0(PC_plus4Reg[28]), .C1(n2131), .Y(n3092) );
  AOI222XL U3354 ( .A0(read_data1[29]), .A1(n2132), .B0(PC_plus4[29]), .B1(
        n3035), .C0(PC_plus4Reg[29]), .C1(n2131), .Y(n3094) );
  AOI222XL U3355 ( .A0(read_data1[30]), .A1(n2132), .B0(PC_plus4[30]), .B1(
        n3035), .C0(PC_plus4Reg[30]), .C1(n2131), .Y(n3096) );
  OAI211X1 U3356 ( .A0(n3220), .A1(n2139), .B0(n3097), .C0(n3098), .Y(n1323)
         );
  AOI222XL U3357 ( .A0(read_data1[31]), .A1(n2132), .B0(PC_plus4[31]), .B1(
        n3035), .C0(PC_plus4Reg[31]), .C1(n2131), .Y(n3098) );
  CLKINVX1 U3358 ( .A(Jump[0]), .Y(n3099) );
  OAI21XL U3359 ( .A0(Jump[1]), .A1(Jump[0]), .B0(n2140), .Y(n3100) );
  NAND2X1 U3360 ( .A(BranchAddr[31]), .B(n3036), .Y(n3097) );
  NOR3X1 U3361 ( .A(WB_Rd[1]), .B(WB_Rd[2]), .C(WB_Rd[0]), .Y(n3002) );
  CLKINVX1 U3362 ( .A(WB_Rd[1]), .Y(n3110) );
  CLKINVX1 U3363 ( .A(WB_Rd[2]), .Y(n3107) );
  CLKINVX1 U3364 ( .A(WB_Rd[0]), .Y(n3109) );
  CLKINVX1 U3365 ( .A(WB_Rd[3]), .Y(n3015) );
  NAND2BX1 U3366 ( .AN(Foward_A[1]), .B(Foward_A[0]), .Y(n3120) );
  NAND2BX1 U3367 ( .AN(Foward_A[0]), .B(Foward_A[1]), .Y(n3118) );
  OAI21XL U3368 ( .A0(n2208), .A1(n3117), .B0(n3184), .Y(after_B_mux[9]) );
  AOI222XL U3369 ( .A0(WB_ALUOut[9]), .A1(n3186), .B0(WB_readdata[9]), .B1(
        n2207), .C0(WB_pcplus4[9]), .C1(n2205), .Y(n2927) );
  CLKMX2X2 U3370 ( .A(after_B_mux[8]), .B(EX_signextend[8]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[8]) );
  OAI21XL U3371 ( .A0(n2208), .A1(n3121), .B0(n3189), .Y(after_B_mux[8]) );
  AOI222XL U3372 ( .A0(WB_ALUOut[8]), .A1(n3186), .B0(WB_readdata[8]), .B1(
        n2207), .C0(WB_pcplus4[8]), .C1(n2205), .Y(n2929) );
  CLKMX2X2 U3373 ( .A(after_B_mux[7]), .B(EX_signextend[7]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[7]) );
  OAI21XL U3374 ( .A0(n2208), .A1(n3123), .B0(n3190), .Y(after_B_mux[7]) );
  AOI222XL U3375 ( .A0(WB_ALUOut[7]), .A1(n3186), .B0(WB_readdata[7]), .B1(
        n2207), .C0(WB_pcplus4[7]), .C1(n2205), .Y(n2930) );
  CLKMX2X2 U3376 ( .A(after_B_mux[6]), .B(EX_signextend[6]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[6]) );
  OAI21XL U3377 ( .A0(n2208), .A1(n3125), .B0(n3191), .Y(after_B_mux[6]) );
  AOI222XL U3378 ( .A0(WB_ALUOut[6]), .A1(n3186), .B0(WB_readdata[6]), .B1(
        n2207), .C0(WB_pcplus4[6]), .C1(n2205), .Y(n2931) );
  CLKINVX1 U3379 ( .A(DCACHE_addr[4]), .Y(n3125) );
  OAI21XL U3380 ( .A0(n2208), .A1(n3127), .B0(n3192), .Y(after_B_mux[5]) );
  AOI222XL U3381 ( .A0(WB_ALUOut[5]), .A1(n3186), .B0(WB_readdata[5]), .B1(
        n2207), .C0(WB_pcplus4[5]), .C1(n2205), .Y(n2932) );
  CLKINVX1 U3382 ( .A(DCACHE_addr[3]), .Y(n3127) );
  OAI21XL U3383 ( .A0(n2208), .A1(n3129), .B0(n3193), .Y(after_B_mux[4]) );
  AOI222XL U3384 ( .A0(WB_ALUOut[4]), .A1(n3186), .B0(WB_readdata[4]), .B1(
        n2207), .C0(WB_pcplus4[4]), .C1(n2205), .Y(n2933) );
  CLKINVX1 U3385 ( .A(DCACHE_addr[2]), .Y(n3129) );
  OAI21XL U3386 ( .A0(n2208), .A1(n3131), .B0(n3194), .Y(after_B_mux[3]) );
  AOI222XL U3387 ( .A0(WB_ALUOut[3]), .A1(n3186), .B0(WB_readdata[3]), .B1(
        n2207), .C0(WB_pcplus4[3]), .C1(n2205), .Y(n2934) );
  CLKMX2X2 U3388 ( .A(after_B_mux[31]), .B(EX_signextend[31]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[31]) );
  OAI21XL U3389 ( .A0(n2208), .A1(n3133), .B0(n3195), .Y(after_B_mux[31]) );
  AOI222XL U3390 ( .A0(WB_ALUOut[31]), .A1(n3186), .B0(WB_readdata[31]), .B1(
        n2207), .C0(WB_pcplus4[31]), .C1(n2205), .Y(n2935) );
  CLKMX2X2 U3391 ( .A(after_B_mux[30]), .B(EX_signextend[30]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[30]) );
  OAI21XL U3392 ( .A0(n2208), .A1(n3135), .B0(n3196), .Y(after_B_mux[30]) );
  AOI222XL U3393 ( .A0(WB_ALUOut[30]), .A1(n3186), .B0(WB_readdata[30]), .B1(
        n2207), .C0(WB_pcplus4[30]), .C1(n2205), .Y(n2936) );
  OAI21XL U3394 ( .A0(n2208), .A1(n3137), .B0(n3197), .Y(after_B_mux[2]) );
  AOI222XL U3395 ( .A0(WB_ALUOut[2]), .A1(n3186), .B0(WB_readdata[2]), .B1(
        n2207), .C0(WB_pcplus4[2]), .C1(n2205), .Y(n2937) );
  OAI21XL U3396 ( .A0(n2208), .A1(n3139), .B0(n3198), .Y(after_B_mux[29]) );
  AOI222XL U3397 ( .A0(WB_ALUOut[29]), .A1(n3186), .B0(WB_readdata[29]), .B1(
        n2207), .C0(WB_pcplus4[29]), .C1(n2205), .Y(n2938) );
  OAI21XL U3398 ( .A0(n2208), .A1(n3141), .B0(n3199), .Y(after_B_mux[28]) );
  AOI222XL U3399 ( .A0(WB_ALUOut[28]), .A1(n3186), .B0(WB_readdata[28]), .B1(
        n2207), .C0(WB_pcplus4[28]), .C1(n2205), .Y(n2939) );
  OAI21XL U3400 ( .A0(n2208), .A1(n3143), .B0(n3200), .Y(after_B_mux[27]) );
  AOI222XL U3401 ( .A0(WB_ALUOut[27]), .A1(n3186), .B0(WB_readdata[27]), .B1(
        n2207), .C0(WB_pcplus4[27]), .C1(n2205), .Y(n2940) );
  OAI21XL U3402 ( .A0(n2208), .A1(n3145), .B0(n3201), .Y(after_B_mux[26]) );
  AOI222XL U3403 ( .A0(WB_ALUOut[26]), .A1(n3186), .B0(WB_readdata[26]), .B1(
        n2207), .C0(WB_pcplus4[26]), .C1(n2205), .Y(n2941) );
  CLKMX2X2 U3404 ( .A(after_B_mux[25]), .B(EX_signextend[25]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[25]) );
  OAI21XL U3405 ( .A0(n2208), .A1(n3147), .B0(n3202), .Y(after_B_mux[25]) );
  AOI222XL U3406 ( .A0(WB_ALUOut[25]), .A1(n3186), .B0(WB_readdata[25]), .B1(
        n2207), .C0(WB_pcplus4[25]), .C1(n2205), .Y(n2942) );
  CLKMX2X2 U3407 ( .A(after_B_mux[24]), .B(EX_signextend[24]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[24]) );
  OAI21XL U3408 ( .A0(n2208), .A1(n3149), .B0(n3203), .Y(after_B_mux[24]) );
  AOI222XL U3409 ( .A0(WB_ALUOut[24]), .A1(n3186), .B0(WB_readdata[24]), .B1(
        n2207), .C0(WB_pcplus4[24]), .C1(n2205), .Y(n2943) );
  CLKMX2X2 U3410 ( .A(after_B_mux[23]), .B(EX_signextend[23]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[23]) );
  OAI21XL U3411 ( .A0(n2208), .A1(n3151), .B0(n3204), .Y(after_B_mux[23]) );
  AOI222XL U3412 ( .A0(WB_ALUOut[23]), .A1(n3186), .B0(WB_readdata[23]), .B1(
        n2207), .C0(WB_pcplus4[23]), .C1(n2205), .Y(n2944) );
  CLKMX2X2 U3413 ( .A(after_B_mux[22]), .B(EX_signextend[22]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[22]) );
  OAI21XL U3414 ( .A0(n2208), .A1(n3153), .B0(n3205), .Y(after_B_mux[22]) );
  AOI222XL U3415 ( .A0(WB_ALUOut[22]), .A1(n3186), .B0(WB_readdata[22]), .B1(
        n2207), .C0(WB_pcplus4[22]), .C1(n2205), .Y(n2945) );
  OAI21XL U3416 ( .A0(n2208), .A1(n3155), .B0(n3206), .Y(after_B_mux[21]) );
  AOI222XL U3417 ( .A0(WB_ALUOut[21]), .A1(n3186), .B0(WB_readdata[21]), .B1(
        n2207), .C0(WB_pcplus4[21]), .C1(n2205), .Y(n2946) );
  OAI21XL U3418 ( .A0(n2208), .A1(n3157), .B0(n3207), .Y(after_B_mux[20]) );
  AOI222XL U3419 ( .A0(WB_ALUOut[20]), .A1(n3186), .B0(WB_readdata[20]), .B1(
        n2207), .C0(WB_pcplus4[20]), .C1(n2205), .Y(n2947) );
  OAI21XL U3420 ( .A0(n2208), .A1(n3159), .B0(n3208), .Y(after_B_mux[1]) );
  AOI222XL U3421 ( .A0(WB_ALUOut[1]), .A1(n3186), .B0(WB_readdata[1]), .B1(
        n2207), .C0(WB_pcplus4[1]), .C1(n2205), .Y(n2948) );
  CLKINVX1 U3422 ( .A(ALUOut_reg[1]), .Y(n3159) );
  OAI21XL U3423 ( .A0(n2208), .A1(n3161), .B0(n3209), .Y(after_B_mux[19]) );
  AOI222XL U3424 ( .A0(WB_ALUOut[19]), .A1(n3186), .B0(WB_readdata[19]), .B1(
        n2207), .C0(WB_pcplus4[19]), .C1(n2205), .Y(n2949) );
  CLKMX2X2 U3425 ( .A(after_B_mux[18]), .B(EX_signextend[18]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[18]) );
  OAI21XL U3426 ( .A0(n2208), .A1(n3163), .B0(n3210), .Y(after_B_mux[18]) );
  AOI222XL U3427 ( .A0(WB_ALUOut[18]), .A1(n3186), .B0(WB_readdata[18]), .B1(
        n2207), .C0(WB_pcplus4[18]), .C1(n2205), .Y(n2950) );
  CLKMX2X2 U3428 ( .A(after_B_mux[17]), .B(EX_signextend[17]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[17]) );
  OAI21XL U3429 ( .A0(n2208), .A1(n3165), .B0(n3211), .Y(after_B_mux[17]) );
  AOI222XL U3430 ( .A0(WB_ALUOut[17]), .A1(n3186), .B0(WB_readdata[17]), .B1(
        n2207), .C0(WB_pcplus4[17]), .C1(n2205), .Y(n2951) );
  CLKMX2X2 U3431 ( .A(after_B_mux[16]), .B(EX_signextend[16]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[16]) );
  OAI21XL U3432 ( .A0(n2208), .A1(n3167), .B0(n3212), .Y(after_B_mux[16]) );
  AOI222XL U3433 ( .A0(WB_ALUOut[16]), .A1(n3186), .B0(WB_readdata[16]), .B1(
        n2207), .C0(WB_pcplus4[16]), .C1(n2205), .Y(n2952) );
  CLKMX2X2 U3434 ( .A(after_B_mux[15]), .B(EX_signextend[15]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[15]) );
  OAI21XL U3435 ( .A0(n2208), .A1(n3169), .B0(n3213), .Y(after_B_mux[15]) );
  AOI222XL U3436 ( .A0(WB_ALUOut[15]), .A1(n3186), .B0(WB_readdata[15]), .B1(
        n2207), .C0(WB_pcplus4[15]), .C1(n2205), .Y(n2953) );
  CLKMX2X2 U3437 ( .A(after_B_mux[14]), .B(EX_signextend[14]), .S0(EX_reg[3]), 
        .Y(after_ALUSrc[14]) );
  OAI21XL U3438 ( .A0(n2208), .A1(n3171), .B0(n3214), .Y(after_B_mux[14]) );
  AOI222XL U3439 ( .A0(WB_ALUOut[14]), .A1(n3186), .B0(WB_readdata[14]), .B1(
        n2207), .C0(WB_pcplus4[14]), .C1(n2205), .Y(n2954) );
  OAI21XL U3440 ( .A0(n2208), .A1(n3173), .B0(n3215), .Y(after_B_mux[13]) );
  AOI222XL U3441 ( .A0(WB_ALUOut[13]), .A1(n3186), .B0(WB_readdata[13]), .B1(
        n2207), .C0(WB_pcplus4[13]), .C1(n2205), .Y(n2955) );
  OAI21XL U3442 ( .A0(n2208), .A1(n3175), .B0(n3216), .Y(after_B_mux[12]) );
  AOI222XL U3443 ( .A0(WB_ALUOut[12]), .A1(n3186), .B0(WB_readdata[12]), .B1(
        n2207), .C0(WB_pcplus4[12]), .C1(n2205), .Y(n2956) );
  OAI21XL U3444 ( .A0(n2208), .A1(n3177), .B0(n3217), .Y(after_B_mux[11]) );
  AOI222XL U3445 ( .A0(WB_ALUOut[11]), .A1(n3186), .B0(WB_readdata[11]), .B1(
        n2207), .C0(WB_pcplus4[11]), .C1(n2205), .Y(n2957) );
  OAI21XL U3446 ( .A0(n2208), .A1(n3179), .B0(n3218), .Y(after_B_mux[10]) );
  AOI222XL U3447 ( .A0(WB_ALUOut[10]), .A1(n3186), .B0(WB_readdata[10]), .B1(
        n2207), .C0(WB_pcplus4[10]), .C1(n2205), .Y(n2958) );
  OAI21XL U3448 ( .A0(n2208), .A1(n3181), .B0(n3219), .Y(after_B_mux[0]) );
  NAND2BX1 U3449 ( .AN(Foward_B[1]), .B(Foward_B[0]), .Y(n3185) );
  AOI222XL U3450 ( .A0(WB_ALUOut[0]), .A1(n3186), .B0(WB_readdata[0]), .B1(
        n2207), .C0(WB_pcplus4[0]), .C1(n2205), .Y(n2959) );
  NOR2BX1 U3451 ( .AN(WB_WB[2]), .B(WB_WB[1]), .Y(n3188) );
  NOR2BX1 U3452 ( .AN(WB_WB[1]), .B(WB_WB[2]), .Y(n3187) );
  CLKINVX1 U3453 ( .A(ALUOut_reg[0]), .Y(n3181) );
  NAND2BX1 U3454 ( .AN(Foward_B[0]), .B(Foward_B[1]), .Y(n3183) );
  AND2X1 U3455 ( .A(M[0]), .B(PCWrite), .Y(MEM_after_detect[0]) );
  AND2X1 U3456 ( .A(RegDST[1]), .B(PCWrite), .Y(WB_after_detect[2]) );
endmodule


module cache_0 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N30, N31, N32, n3804, \CACHE[7][154] , \CACHE[7][153] ,
         \CACHE[7][152] , \CACHE[7][151] , \CACHE[7][150] , \CACHE[7][149] ,
         \CACHE[7][148] , \CACHE[7][147] , \CACHE[7][146] , \CACHE[7][145] ,
         \CACHE[7][144] , \CACHE[7][143] , \CACHE[7][142] , \CACHE[7][141] ,
         \CACHE[7][140] , \CACHE[7][139] , \CACHE[7][138] , \CACHE[7][137] ,
         \CACHE[7][136] , \CACHE[7][135] , \CACHE[7][134] , \CACHE[7][133] ,
         \CACHE[7][132] , \CACHE[7][131] , \CACHE[7][130] , \CACHE[7][129] ,
         \CACHE[7][128] , \CACHE[7][127] , \CACHE[7][126] , \CACHE[7][125] ,
         \CACHE[7][124] , \CACHE[7][123] , \CACHE[7][122] , \CACHE[7][121] ,
         \CACHE[7][120] , \CACHE[7][119] , \CACHE[7][118] , \CACHE[7][117] ,
         \CACHE[7][116] , \CACHE[7][115] , \CACHE[7][114] , \CACHE[7][113] ,
         \CACHE[7][112] , \CACHE[7][111] , \CACHE[7][110] , \CACHE[7][109] ,
         \CACHE[7][108] , \CACHE[7][107] , \CACHE[7][106] , \CACHE[7][105] ,
         \CACHE[7][104] , \CACHE[7][103] , \CACHE[7][102] , \CACHE[7][101] ,
         \CACHE[7][100] , \CACHE[7][99] , \CACHE[7][98] , \CACHE[7][97] ,
         \CACHE[7][96] , \CACHE[7][95] , \CACHE[7][94] , \CACHE[7][93] ,
         \CACHE[7][92] , \CACHE[7][91] , \CACHE[7][90] , \CACHE[7][89] ,
         \CACHE[7][88] , \CACHE[7][87] , \CACHE[7][86] , \CACHE[7][85] ,
         \CACHE[7][84] , \CACHE[7][83] , \CACHE[7][82] , \CACHE[7][81] ,
         \CACHE[7][80] , \CACHE[7][79] , \CACHE[7][78] , \CACHE[7][77] ,
         \CACHE[7][76] , \CACHE[7][75] , \CACHE[7][74] , \CACHE[7][73] ,
         \CACHE[7][72] , \CACHE[7][71] , \CACHE[7][70] , \CACHE[7][69] ,
         \CACHE[7][68] , \CACHE[7][67] , \CACHE[7][66] , \CACHE[7][65] ,
         \CACHE[7][64] , \CACHE[7][63] , \CACHE[7][62] , \CACHE[7][61] ,
         \CACHE[7][60] , \CACHE[7][59] , \CACHE[7][58] , \CACHE[7][57] ,
         \CACHE[7][56] , \CACHE[7][55] , \CACHE[7][54] , \CACHE[7][53] ,
         \CACHE[7][52] , \CACHE[7][51] , \CACHE[7][50] , \CACHE[7][49] ,
         \CACHE[7][48] , \CACHE[7][47] , \CACHE[7][46] , \CACHE[7][45] ,
         \CACHE[7][44] , \CACHE[7][43] , \CACHE[7][42] , \CACHE[7][41] ,
         \CACHE[7][40] , \CACHE[7][39] , \CACHE[7][38] , \CACHE[7][37] ,
         \CACHE[7][36] , \CACHE[7][35] , \CACHE[7][34] , \CACHE[7][33] ,
         \CACHE[7][32] , \CACHE[7][31] , \CACHE[7][30] , \CACHE[7][29] ,
         \CACHE[7][28] , \CACHE[7][27] , \CACHE[7][26] , \CACHE[7][25] ,
         \CACHE[7][24] , \CACHE[7][23] , \CACHE[7][22] , \CACHE[7][21] ,
         \CACHE[7][20] , \CACHE[7][19] , \CACHE[7][18] , \CACHE[7][17] ,
         \CACHE[7][16] , \CACHE[7][15] , \CACHE[7][14] , \CACHE[7][13] ,
         \CACHE[7][12] , \CACHE[7][11] , \CACHE[7][10] , \CACHE[7][9] ,
         \CACHE[7][8] , \CACHE[7][7] , \CACHE[7][6] , \CACHE[7][5] ,
         \CACHE[7][4] , \CACHE[7][3] , \CACHE[7][2] , \CACHE[7][1] ,
         \CACHE[7][0] , \CACHE[6][154] , \CACHE[6][153] , \CACHE[6][152] ,
         \CACHE[6][151] , \CACHE[6][150] , \CACHE[6][149] , \CACHE[6][148] ,
         \CACHE[6][147] , \CACHE[6][146] , \CACHE[6][145] , \CACHE[6][144] ,
         \CACHE[6][143] , \CACHE[6][142] , \CACHE[6][141] , \CACHE[6][140] ,
         \CACHE[6][139] , \CACHE[6][138] , \CACHE[6][137] , \CACHE[6][136] ,
         \CACHE[6][135] , \CACHE[6][134] , \CACHE[6][133] , \CACHE[6][132] ,
         \CACHE[6][131] , \CACHE[6][130] , \CACHE[6][129] , \CACHE[6][128] ,
         \CACHE[6][127] , \CACHE[6][126] , \CACHE[6][125] , \CACHE[6][124] ,
         \CACHE[6][123] , \CACHE[6][122] , \CACHE[6][121] , \CACHE[6][120] ,
         \CACHE[6][119] , \CACHE[6][118] , \CACHE[6][117] , \CACHE[6][116] ,
         \CACHE[6][115] , \CACHE[6][114] , \CACHE[6][113] , \CACHE[6][112] ,
         \CACHE[6][111] , \CACHE[6][110] , \CACHE[6][109] , \CACHE[6][108] ,
         \CACHE[6][107] , \CACHE[6][106] , \CACHE[6][105] , \CACHE[6][104] ,
         \CACHE[6][103] , \CACHE[6][102] , \CACHE[6][101] , \CACHE[6][100] ,
         \CACHE[6][99] , \CACHE[6][98] , \CACHE[6][97] , \CACHE[6][96] ,
         \CACHE[6][95] , \CACHE[6][94] , \CACHE[6][93] , \CACHE[6][92] ,
         \CACHE[6][91] , \CACHE[6][90] , \CACHE[6][89] , \CACHE[6][88] ,
         \CACHE[6][87] , \CACHE[6][86] , \CACHE[6][85] , \CACHE[6][84] ,
         \CACHE[6][83] , \CACHE[6][82] , \CACHE[6][81] , \CACHE[6][80] ,
         \CACHE[6][79] , \CACHE[6][78] , \CACHE[6][77] , \CACHE[6][76] ,
         \CACHE[6][75] , \CACHE[6][74] , \CACHE[6][73] , \CACHE[6][72] ,
         \CACHE[6][71] , \CACHE[6][70] , \CACHE[6][69] , \CACHE[6][68] ,
         \CACHE[6][67] , \CACHE[6][66] , \CACHE[6][65] , \CACHE[6][64] ,
         \CACHE[6][63] , \CACHE[6][62] , \CACHE[6][61] , \CACHE[6][60] ,
         \CACHE[6][59] , \CACHE[6][58] , \CACHE[6][57] , \CACHE[6][56] ,
         \CACHE[6][55] , \CACHE[6][54] , \CACHE[6][53] , \CACHE[6][52] ,
         \CACHE[6][51] , \CACHE[6][50] , \CACHE[6][49] , \CACHE[6][48] ,
         \CACHE[6][47] , \CACHE[6][46] , \CACHE[6][45] , \CACHE[6][44] ,
         \CACHE[6][43] , \CACHE[6][42] , \CACHE[6][41] , \CACHE[6][40] ,
         \CACHE[6][39] , \CACHE[6][38] , \CACHE[6][37] , \CACHE[6][36] ,
         \CACHE[6][35] , \CACHE[6][34] , \CACHE[6][33] , \CACHE[6][32] ,
         \CACHE[6][31] , \CACHE[6][30] , \CACHE[6][29] , \CACHE[6][28] ,
         \CACHE[6][27] , \CACHE[6][26] , \CACHE[6][25] , \CACHE[6][24] ,
         \CACHE[6][23] , \CACHE[6][22] , \CACHE[6][21] , \CACHE[6][20] ,
         \CACHE[6][19] , \CACHE[6][18] , \CACHE[6][17] , \CACHE[6][16] ,
         \CACHE[6][15] , \CACHE[6][14] , \CACHE[6][13] , \CACHE[6][12] ,
         \CACHE[6][11] , \CACHE[6][10] , \CACHE[6][9] , \CACHE[6][8] ,
         \CACHE[6][7] , \CACHE[6][6] , \CACHE[6][5] , \CACHE[6][4] ,
         \CACHE[6][3] , \CACHE[6][2] , \CACHE[6][1] , \CACHE[6][0] ,
         \CACHE[5][154] , \CACHE[5][153] , \CACHE[5][152] , \CACHE[5][151] ,
         \CACHE[5][150] , \CACHE[5][149] , \CACHE[5][148] , \CACHE[5][147] ,
         \CACHE[5][146] , \CACHE[5][145] , \CACHE[5][144] , \CACHE[5][143] ,
         \CACHE[5][142] , \CACHE[5][141] , \CACHE[5][140] , \CACHE[5][139] ,
         \CACHE[5][138] , \CACHE[5][137] , \CACHE[5][136] , \CACHE[5][135] ,
         \CACHE[5][134] , \CACHE[5][133] , \CACHE[5][132] , \CACHE[5][131] ,
         \CACHE[5][130] , \CACHE[5][129] , \CACHE[5][128] , \CACHE[5][127] ,
         \CACHE[5][126] , \CACHE[5][125] , \CACHE[5][124] , \CACHE[5][123] ,
         \CACHE[5][122] , \CACHE[5][121] , \CACHE[5][120] , \CACHE[5][119] ,
         \CACHE[5][118] , \CACHE[5][117] , \CACHE[5][116] , \CACHE[5][115] ,
         \CACHE[5][114] , \CACHE[5][113] , \CACHE[5][112] , \CACHE[5][111] ,
         \CACHE[5][110] , \CACHE[5][109] , \CACHE[5][108] , \CACHE[5][107] ,
         \CACHE[5][106] , \CACHE[5][105] , \CACHE[5][104] , \CACHE[5][103] ,
         \CACHE[5][102] , \CACHE[5][101] , \CACHE[5][100] , \CACHE[5][99] ,
         \CACHE[5][98] , \CACHE[5][97] , \CACHE[5][96] , \CACHE[5][95] ,
         \CACHE[5][94] , \CACHE[5][93] , \CACHE[5][92] , \CACHE[5][91] ,
         \CACHE[5][90] , \CACHE[5][89] , \CACHE[5][88] , \CACHE[5][87] ,
         \CACHE[5][86] , \CACHE[5][85] , \CACHE[5][84] , \CACHE[5][83] ,
         \CACHE[5][82] , \CACHE[5][81] , \CACHE[5][80] , \CACHE[5][79] ,
         \CACHE[5][78] , \CACHE[5][77] , \CACHE[5][76] , \CACHE[5][75] ,
         \CACHE[5][74] , \CACHE[5][73] , \CACHE[5][72] , \CACHE[5][71] ,
         \CACHE[5][70] , \CACHE[5][69] , \CACHE[5][68] , \CACHE[5][67] ,
         \CACHE[5][66] , \CACHE[5][65] , \CACHE[5][64] , \CACHE[5][63] ,
         \CACHE[5][62] , \CACHE[5][61] , \CACHE[5][60] , \CACHE[5][59] ,
         \CACHE[5][58] , \CACHE[5][57] , \CACHE[5][56] , \CACHE[5][55] ,
         \CACHE[5][54] , \CACHE[5][53] , \CACHE[5][52] , \CACHE[5][51] ,
         \CACHE[5][50] , \CACHE[5][49] , \CACHE[5][48] , \CACHE[5][47] ,
         \CACHE[5][46] , \CACHE[5][45] , \CACHE[5][44] , \CACHE[5][43] ,
         \CACHE[5][42] , \CACHE[5][41] , \CACHE[5][40] , \CACHE[5][39] ,
         \CACHE[5][38] , \CACHE[5][37] , \CACHE[5][36] , \CACHE[5][35] ,
         \CACHE[5][34] , \CACHE[5][33] , \CACHE[5][32] , \CACHE[5][31] ,
         \CACHE[5][30] , \CACHE[5][29] , \CACHE[5][28] , \CACHE[5][27] ,
         \CACHE[5][26] , \CACHE[5][25] , \CACHE[5][24] , \CACHE[5][23] ,
         \CACHE[5][22] , \CACHE[5][21] , \CACHE[5][20] , \CACHE[5][19] ,
         \CACHE[5][18] , \CACHE[5][17] , \CACHE[5][16] , \CACHE[5][15] ,
         \CACHE[5][14] , \CACHE[5][13] , \CACHE[5][12] , \CACHE[5][11] ,
         \CACHE[5][10] , \CACHE[5][9] , \CACHE[5][8] , \CACHE[5][7] ,
         \CACHE[5][6] , \CACHE[5][5] , \CACHE[5][4] , \CACHE[5][3] ,
         \CACHE[5][2] , \CACHE[5][1] , \CACHE[5][0] , \CACHE[4][154] ,
         \CACHE[4][153] , \CACHE[4][152] , \CACHE[4][151] , \CACHE[4][150] ,
         \CACHE[4][149] , \CACHE[4][148] , \CACHE[4][147] , \CACHE[4][146] ,
         \CACHE[4][145] , \CACHE[4][144] , \CACHE[4][143] , \CACHE[4][142] ,
         \CACHE[4][141] , \CACHE[4][140] , \CACHE[4][139] , \CACHE[4][138] ,
         \CACHE[4][137] , \CACHE[4][136] , \CACHE[4][135] , \CACHE[4][134] ,
         \CACHE[4][133] , \CACHE[4][132] , \CACHE[4][131] , \CACHE[4][130] ,
         \CACHE[4][129] , \CACHE[4][128] , \CACHE[4][127] , \CACHE[4][126] ,
         \CACHE[4][125] , \CACHE[4][124] , \CACHE[4][123] , \CACHE[4][122] ,
         \CACHE[4][121] , \CACHE[4][120] , \CACHE[4][119] , \CACHE[4][118] ,
         \CACHE[4][117] , \CACHE[4][116] , \CACHE[4][115] , \CACHE[4][114] ,
         \CACHE[4][113] , \CACHE[4][112] , \CACHE[4][111] , \CACHE[4][110] ,
         \CACHE[4][109] , \CACHE[4][108] , \CACHE[4][107] , \CACHE[4][106] ,
         \CACHE[4][105] , \CACHE[4][104] , \CACHE[4][103] , \CACHE[4][102] ,
         \CACHE[4][101] , \CACHE[4][100] , \CACHE[4][99] , \CACHE[4][98] ,
         \CACHE[4][97] , \CACHE[4][96] , \CACHE[4][95] , \CACHE[4][94] ,
         \CACHE[4][93] , \CACHE[4][92] , \CACHE[4][91] , \CACHE[4][90] ,
         \CACHE[4][89] , \CACHE[4][88] , \CACHE[4][87] , \CACHE[4][86] ,
         \CACHE[4][85] , \CACHE[4][84] , \CACHE[4][83] , \CACHE[4][82] ,
         \CACHE[4][81] , \CACHE[4][80] , \CACHE[4][79] , \CACHE[4][78] ,
         \CACHE[4][77] , \CACHE[4][76] , \CACHE[4][75] , \CACHE[4][74] ,
         \CACHE[4][73] , \CACHE[4][72] , \CACHE[4][71] , \CACHE[4][70] ,
         \CACHE[4][69] , \CACHE[4][68] , \CACHE[4][67] , \CACHE[4][66] ,
         \CACHE[4][65] , \CACHE[4][64] , \CACHE[4][63] , \CACHE[4][62] ,
         \CACHE[4][61] , \CACHE[4][60] , \CACHE[4][59] , \CACHE[4][58] ,
         \CACHE[4][57] , \CACHE[4][56] , \CACHE[4][55] , \CACHE[4][54] ,
         \CACHE[4][53] , \CACHE[4][52] , \CACHE[4][51] , \CACHE[4][50] ,
         \CACHE[4][49] , \CACHE[4][48] , \CACHE[4][47] , \CACHE[4][46] ,
         \CACHE[4][45] , \CACHE[4][44] , \CACHE[4][43] , \CACHE[4][42] ,
         \CACHE[4][41] , \CACHE[4][40] , \CACHE[4][39] , \CACHE[4][38] ,
         \CACHE[4][37] , \CACHE[4][36] , \CACHE[4][35] , \CACHE[4][34] ,
         \CACHE[4][33] , \CACHE[4][32] , \CACHE[4][31] , \CACHE[4][30] ,
         \CACHE[4][29] , \CACHE[4][28] , \CACHE[4][27] , \CACHE[4][26] ,
         \CACHE[4][25] , \CACHE[4][24] , \CACHE[4][23] , \CACHE[4][22] ,
         \CACHE[4][21] , \CACHE[4][20] , \CACHE[4][19] , \CACHE[4][18] ,
         \CACHE[4][17] , \CACHE[4][16] , \CACHE[4][15] , \CACHE[4][14] ,
         \CACHE[4][13] , \CACHE[4][12] , \CACHE[4][11] , \CACHE[4][10] ,
         \CACHE[4][9] , \CACHE[4][8] , \CACHE[4][7] , \CACHE[4][6] ,
         \CACHE[4][5] , \CACHE[4][4] , \CACHE[4][3] , \CACHE[4][2] ,
         \CACHE[4][1] , \CACHE[4][0] , \CACHE[3][154] , \CACHE[3][153] ,
         \CACHE[3][152] , \CACHE[3][151] , \CACHE[3][150] , \CACHE[3][149] ,
         \CACHE[3][148] , \CACHE[3][147] , \CACHE[3][146] , \CACHE[3][145] ,
         \CACHE[3][144] , \CACHE[3][143] , \CACHE[3][142] , \CACHE[3][141] ,
         \CACHE[3][140] , \CACHE[3][139] , \CACHE[3][138] , \CACHE[3][137] ,
         \CACHE[3][136] , \CACHE[3][135] , \CACHE[3][134] , \CACHE[3][133] ,
         \CACHE[3][132] , \CACHE[3][131] , \CACHE[3][130] , \CACHE[3][129] ,
         \CACHE[3][128] , \CACHE[3][127] , \CACHE[3][126] , \CACHE[3][125] ,
         \CACHE[3][124] , \CACHE[3][123] , \CACHE[3][122] , \CACHE[3][121] ,
         \CACHE[3][120] , \CACHE[3][119] , \CACHE[3][118] , \CACHE[3][117] ,
         \CACHE[3][116] , \CACHE[3][115] , \CACHE[3][114] , \CACHE[3][113] ,
         \CACHE[3][112] , \CACHE[3][111] , \CACHE[3][110] , \CACHE[3][109] ,
         \CACHE[3][108] , \CACHE[3][107] , \CACHE[3][106] , \CACHE[3][105] ,
         \CACHE[3][104] , \CACHE[3][103] , \CACHE[3][102] , \CACHE[3][101] ,
         \CACHE[3][100] , \CACHE[3][99] , \CACHE[3][98] , \CACHE[3][97] ,
         \CACHE[3][96] , \CACHE[3][95] , \CACHE[3][94] , \CACHE[3][93] ,
         \CACHE[3][92] , \CACHE[3][91] , \CACHE[3][90] , \CACHE[3][89] ,
         \CACHE[3][88] , \CACHE[3][87] , \CACHE[3][86] , \CACHE[3][85] ,
         \CACHE[3][84] , \CACHE[3][83] , \CACHE[3][82] , \CACHE[3][81] ,
         \CACHE[3][80] , \CACHE[3][79] , \CACHE[3][78] , \CACHE[3][77] ,
         \CACHE[3][76] , \CACHE[3][75] , \CACHE[3][74] , \CACHE[3][73] ,
         \CACHE[3][72] , \CACHE[3][71] , \CACHE[3][70] , \CACHE[3][69] ,
         \CACHE[3][68] , \CACHE[3][67] , \CACHE[3][66] , \CACHE[3][65] ,
         \CACHE[3][64] , \CACHE[3][63] , \CACHE[3][62] , \CACHE[3][61] ,
         \CACHE[3][60] , \CACHE[3][59] , \CACHE[3][58] , \CACHE[3][57] ,
         \CACHE[3][56] , \CACHE[3][55] , \CACHE[3][54] , \CACHE[3][53] ,
         \CACHE[3][52] , \CACHE[3][51] , \CACHE[3][50] , \CACHE[3][49] ,
         \CACHE[3][48] , \CACHE[3][47] , \CACHE[3][46] , \CACHE[3][45] ,
         \CACHE[3][44] , \CACHE[3][43] , \CACHE[3][42] , \CACHE[3][41] ,
         \CACHE[3][40] , \CACHE[3][39] , \CACHE[3][38] , \CACHE[3][37] ,
         \CACHE[3][36] , \CACHE[3][35] , \CACHE[3][34] , \CACHE[3][33] ,
         \CACHE[3][32] , \CACHE[3][31] , \CACHE[3][30] , \CACHE[3][29] ,
         \CACHE[3][28] , \CACHE[3][27] , \CACHE[3][26] , \CACHE[3][25] ,
         \CACHE[3][24] , \CACHE[3][23] , \CACHE[3][22] , \CACHE[3][21] ,
         \CACHE[3][20] , \CACHE[3][19] , \CACHE[3][18] , \CACHE[3][17] ,
         \CACHE[3][16] , \CACHE[3][15] , \CACHE[3][14] , \CACHE[3][13] ,
         \CACHE[3][12] , \CACHE[3][11] , \CACHE[3][10] , \CACHE[3][9] ,
         \CACHE[3][8] , \CACHE[3][7] , \CACHE[3][6] , \CACHE[3][5] ,
         \CACHE[3][4] , \CACHE[3][3] , \CACHE[3][2] , \CACHE[3][1] ,
         \CACHE[3][0] , \CACHE[2][154] , \CACHE[2][153] , \CACHE[2][152] ,
         \CACHE[2][151] , \CACHE[2][150] , \CACHE[2][149] , \CACHE[2][148] ,
         \CACHE[2][147] , \CACHE[2][146] , \CACHE[2][145] , \CACHE[2][144] ,
         \CACHE[2][143] , \CACHE[2][142] , \CACHE[2][141] , \CACHE[2][140] ,
         \CACHE[2][139] , \CACHE[2][138] , \CACHE[2][137] , \CACHE[2][136] ,
         \CACHE[2][135] , \CACHE[2][134] , \CACHE[2][133] , \CACHE[2][132] ,
         \CACHE[2][131] , \CACHE[2][130] , \CACHE[2][129] , \CACHE[2][128] ,
         \CACHE[2][127] , \CACHE[2][126] , \CACHE[2][125] , \CACHE[2][124] ,
         \CACHE[2][123] , \CACHE[2][122] , \CACHE[2][121] , \CACHE[2][120] ,
         \CACHE[2][119] , \CACHE[2][118] , \CACHE[2][117] , \CACHE[2][116] ,
         \CACHE[2][115] , \CACHE[2][114] , \CACHE[2][113] , \CACHE[2][112] ,
         \CACHE[2][111] , \CACHE[2][110] , \CACHE[2][109] , \CACHE[2][108] ,
         \CACHE[2][107] , \CACHE[2][106] , \CACHE[2][105] , \CACHE[2][104] ,
         \CACHE[2][103] , \CACHE[2][102] , \CACHE[2][101] , \CACHE[2][100] ,
         \CACHE[2][99] , \CACHE[2][98] , \CACHE[2][97] , \CACHE[2][96] ,
         \CACHE[2][95] , \CACHE[2][94] , \CACHE[2][93] , \CACHE[2][92] ,
         \CACHE[2][91] , \CACHE[2][90] , \CACHE[2][89] , \CACHE[2][88] ,
         \CACHE[2][87] , \CACHE[2][86] , \CACHE[2][85] , \CACHE[2][84] ,
         \CACHE[2][83] , \CACHE[2][82] , \CACHE[2][81] , \CACHE[2][80] ,
         \CACHE[2][79] , \CACHE[2][78] , \CACHE[2][77] , \CACHE[2][76] ,
         \CACHE[2][75] , \CACHE[2][74] , \CACHE[2][73] , \CACHE[2][72] ,
         \CACHE[2][71] , \CACHE[2][70] , \CACHE[2][69] , \CACHE[2][68] ,
         \CACHE[2][67] , \CACHE[2][66] , \CACHE[2][65] , \CACHE[2][64] ,
         \CACHE[2][63] , \CACHE[2][62] , \CACHE[2][61] , \CACHE[2][60] ,
         \CACHE[2][59] , \CACHE[2][58] , \CACHE[2][57] , \CACHE[2][56] ,
         \CACHE[2][55] , \CACHE[2][54] , \CACHE[2][53] , \CACHE[2][52] ,
         \CACHE[2][51] , \CACHE[2][50] , \CACHE[2][49] , \CACHE[2][48] ,
         \CACHE[2][47] , \CACHE[2][46] , \CACHE[2][45] , \CACHE[2][44] ,
         \CACHE[2][43] , \CACHE[2][42] , \CACHE[2][41] , \CACHE[2][40] ,
         \CACHE[2][39] , \CACHE[2][38] , \CACHE[2][37] , \CACHE[2][36] ,
         \CACHE[2][35] , \CACHE[2][34] , \CACHE[2][33] , \CACHE[2][32] ,
         \CACHE[2][31] , \CACHE[2][30] , \CACHE[2][29] , \CACHE[2][28] ,
         \CACHE[2][27] , \CACHE[2][26] , \CACHE[2][25] , \CACHE[2][24] ,
         \CACHE[2][23] , \CACHE[2][22] , \CACHE[2][21] , \CACHE[2][20] ,
         \CACHE[2][19] , \CACHE[2][18] , \CACHE[2][17] , \CACHE[2][16] ,
         \CACHE[2][15] , \CACHE[2][14] , \CACHE[2][13] , \CACHE[2][12] ,
         \CACHE[2][11] , \CACHE[2][10] , \CACHE[2][9] , \CACHE[2][8] ,
         \CACHE[2][7] , \CACHE[2][6] , \CACHE[2][5] , \CACHE[2][4] ,
         \CACHE[2][3] , \CACHE[2][2] , \CACHE[2][1] , \CACHE[2][0] ,
         \CACHE[1][154] , \CACHE[1][153] , \CACHE[1][152] , \CACHE[1][151] ,
         \CACHE[1][150] , \CACHE[1][149] , \CACHE[1][148] , \CACHE[1][147] ,
         \CACHE[1][146] , \CACHE[1][145] , \CACHE[1][144] , \CACHE[1][143] ,
         \CACHE[1][142] , \CACHE[1][141] , \CACHE[1][140] , \CACHE[1][139] ,
         \CACHE[1][138] , \CACHE[1][137] , \CACHE[1][136] , \CACHE[1][135] ,
         \CACHE[1][134] , \CACHE[1][133] , \CACHE[1][132] , \CACHE[1][131] ,
         \CACHE[1][130] , \CACHE[1][129] , \CACHE[1][128] , \CACHE[1][127] ,
         \CACHE[1][126] , \CACHE[1][125] , \CACHE[1][124] , \CACHE[1][123] ,
         \CACHE[1][122] , \CACHE[1][121] , \CACHE[1][120] , \CACHE[1][119] ,
         \CACHE[1][118] , \CACHE[1][117] , \CACHE[1][116] , \CACHE[1][115] ,
         \CACHE[1][114] , \CACHE[1][113] , \CACHE[1][112] , \CACHE[1][111] ,
         \CACHE[1][110] , \CACHE[1][109] , \CACHE[1][108] , \CACHE[1][107] ,
         \CACHE[1][106] , \CACHE[1][105] , \CACHE[1][104] , \CACHE[1][103] ,
         \CACHE[1][102] , \CACHE[1][101] , \CACHE[1][100] , \CACHE[1][99] ,
         \CACHE[1][98] , \CACHE[1][97] , \CACHE[1][96] , \CACHE[1][95] ,
         \CACHE[1][94] , \CACHE[1][93] , \CACHE[1][92] , \CACHE[1][91] ,
         \CACHE[1][90] , \CACHE[1][89] , \CACHE[1][88] , \CACHE[1][87] ,
         \CACHE[1][86] , \CACHE[1][85] , \CACHE[1][84] , \CACHE[1][83] ,
         \CACHE[1][82] , \CACHE[1][81] , \CACHE[1][80] , \CACHE[1][79] ,
         \CACHE[1][78] , \CACHE[1][77] , \CACHE[1][76] , \CACHE[1][75] ,
         \CACHE[1][74] , \CACHE[1][73] , \CACHE[1][72] , \CACHE[1][71] ,
         \CACHE[1][70] , \CACHE[1][69] , \CACHE[1][68] , \CACHE[1][67] ,
         \CACHE[1][66] , \CACHE[1][65] , \CACHE[1][64] , \CACHE[1][63] ,
         \CACHE[1][62] , \CACHE[1][61] , \CACHE[1][60] , \CACHE[1][59] ,
         \CACHE[1][58] , \CACHE[1][57] , \CACHE[1][56] , \CACHE[1][55] ,
         \CACHE[1][54] , \CACHE[1][53] , \CACHE[1][52] , \CACHE[1][51] ,
         \CACHE[1][50] , \CACHE[1][49] , \CACHE[1][48] , \CACHE[1][47] ,
         \CACHE[1][46] , \CACHE[1][45] , \CACHE[1][44] , \CACHE[1][43] ,
         \CACHE[1][42] , \CACHE[1][41] , \CACHE[1][40] , \CACHE[1][39] ,
         \CACHE[1][38] , \CACHE[1][37] , \CACHE[1][36] , \CACHE[1][35] ,
         \CACHE[1][34] , \CACHE[1][33] , \CACHE[1][32] , \CACHE[1][31] ,
         \CACHE[1][30] , \CACHE[1][29] , \CACHE[1][28] , \CACHE[1][27] ,
         \CACHE[1][26] , \CACHE[1][25] , \CACHE[1][24] , \CACHE[1][23] ,
         \CACHE[1][22] , \CACHE[1][21] , \CACHE[1][20] , \CACHE[1][19] ,
         \CACHE[1][18] , \CACHE[1][17] , \CACHE[1][16] , \CACHE[1][15] ,
         \CACHE[1][14] , \CACHE[1][13] , \CACHE[1][12] , \CACHE[1][11] ,
         \CACHE[1][10] , \CACHE[1][9] , \CACHE[1][8] , \CACHE[1][7] ,
         \CACHE[1][6] , \CACHE[1][5] , \CACHE[1][4] , \CACHE[1][3] ,
         \CACHE[1][2] , \CACHE[1][1] , \CACHE[1][0] , \CACHE[0][154] ,
         \CACHE[0][153] , \CACHE[0][152] , \CACHE[0][151] , \CACHE[0][150] ,
         \CACHE[0][149] , \CACHE[0][148] , \CACHE[0][147] , \CACHE[0][146] ,
         \CACHE[0][145] , \CACHE[0][144] , \CACHE[0][143] , \CACHE[0][142] ,
         \CACHE[0][141] , \CACHE[0][140] , \CACHE[0][139] , \CACHE[0][138] ,
         \CACHE[0][137] , \CACHE[0][136] , \CACHE[0][135] , \CACHE[0][134] ,
         \CACHE[0][133] , \CACHE[0][132] , \CACHE[0][131] , \CACHE[0][130] ,
         \CACHE[0][129] , \CACHE[0][128] , \CACHE[0][127] , \CACHE[0][126] ,
         \CACHE[0][125] , \CACHE[0][124] , \CACHE[0][123] , \CACHE[0][122] ,
         \CACHE[0][121] , \CACHE[0][120] , \CACHE[0][119] , \CACHE[0][118] ,
         \CACHE[0][117] , \CACHE[0][116] , \CACHE[0][115] , \CACHE[0][114] ,
         \CACHE[0][113] , \CACHE[0][112] , \CACHE[0][111] , \CACHE[0][110] ,
         \CACHE[0][109] , \CACHE[0][108] , \CACHE[0][107] , \CACHE[0][106] ,
         \CACHE[0][105] , \CACHE[0][104] , \CACHE[0][103] , \CACHE[0][102] ,
         \CACHE[0][101] , \CACHE[0][100] , \CACHE[0][99] , \CACHE[0][98] ,
         \CACHE[0][97] , \CACHE[0][96] , \CACHE[0][95] , \CACHE[0][94] ,
         \CACHE[0][93] , \CACHE[0][92] , \CACHE[0][91] , \CACHE[0][90] ,
         \CACHE[0][89] , \CACHE[0][88] , \CACHE[0][87] , \CACHE[0][86] ,
         \CACHE[0][85] , \CACHE[0][84] , \CACHE[0][83] , \CACHE[0][82] ,
         \CACHE[0][81] , \CACHE[0][80] , \CACHE[0][79] , \CACHE[0][78] ,
         \CACHE[0][77] , \CACHE[0][76] , \CACHE[0][75] , \CACHE[0][74] ,
         \CACHE[0][73] , \CACHE[0][72] , \CACHE[0][71] , \CACHE[0][70] ,
         \CACHE[0][69] , \CACHE[0][68] , \CACHE[0][67] , \CACHE[0][66] ,
         \CACHE[0][65] , \CACHE[0][64] , \CACHE[0][63] , \CACHE[0][62] ,
         \CACHE[0][61] , \CACHE[0][60] , \CACHE[0][59] , \CACHE[0][58] ,
         \CACHE[0][57] , \CACHE[0][56] , \CACHE[0][55] , \CACHE[0][54] ,
         \CACHE[0][53] , \CACHE[0][52] , \CACHE[0][51] , \CACHE[0][50] ,
         \CACHE[0][49] , \CACHE[0][48] , \CACHE[0][47] , \CACHE[0][46] ,
         \CACHE[0][45] , \CACHE[0][44] , \CACHE[0][43] , \CACHE[0][42] ,
         \CACHE[0][41] , \CACHE[0][40] , \CACHE[0][39] , \CACHE[0][38] ,
         \CACHE[0][37] , \CACHE[0][36] , \CACHE[0][35] , \CACHE[0][34] ,
         \CACHE[0][33] , \CACHE[0][32] , \CACHE[0][31] , \CACHE[0][30] ,
         \CACHE[0][29] , \CACHE[0][28] , \CACHE[0][27] , \CACHE[0][26] ,
         \CACHE[0][25] , \CACHE[0][24] , \CACHE[0][23] , \CACHE[0][22] ,
         \CACHE[0][21] , \CACHE[0][20] , \CACHE[0][19] , \CACHE[0][18] ,
         \CACHE[0][17] , \CACHE[0][16] , \CACHE[0][15] , \CACHE[0][14] ,
         \CACHE[0][13] , \CACHE[0][12] , \CACHE[0][11] , \CACHE[0][10] ,
         \CACHE[0][9] , \CACHE[0][8] , \CACHE[0][7] , \CACHE[0][6] ,
         \CACHE[0][5] , \CACHE[0][4] , \CACHE[0][3] , \CACHE[0][2] ,
         \CACHE[0][1] , \CACHE[0][0] , N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96,
         N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108,
         N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119,
         N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130,
         N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141,
         N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152,
         N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163,
         N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174,
         N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185,
         N186, N187, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3021,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n316, n317, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n3020, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803;
  assign N30 = proc_addr[2];
  assign N31 = proc_addr[3];
  assign N32 = proc_addr[4];

  DFFRX1 \CACHE_reg[7][154]  ( .D(n3021), .CK(clk), .RN(n3057), .Q(
        \CACHE[7][154] ), .QN(n1780) );
  DFFRX1 \CACHE_reg[7][153]  ( .D(n3019), .CK(clk), .RN(n3056), .Q(
        \CACHE[7][153] ), .QN(n1779) );
  DFFRX1 \CACHE_reg[7][152]  ( .D(n3018), .CK(clk), .RN(n3056), .Q(
        \CACHE[7][152] ), .QN(n1778) );
  DFFRX1 \CACHE_reg[7][151]  ( .D(n3017), .CK(clk), .RN(n3040), .Q(
        \CACHE[7][151] ), .QN(n1777) );
  DFFRX1 \CACHE_reg[7][150]  ( .D(n3016), .CK(clk), .RN(n3040), .Q(
        \CACHE[7][150] ), .QN(n1776) );
  DFFRX1 \CACHE_reg[7][149]  ( .D(n3015), .CK(clk), .RN(n3041), .Q(
        \CACHE[7][149] ), .QN(n1775) );
  DFFRX1 \CACHE_reg[7][148]  ( .D(n3014), .CK(clk), .RN(n3042), .Q(
        \CACHE[7][148] ), .QN(n1774) );
  DFFRX1 \CACHE_reg[7][147]  ( .D(n3013), .CK(clk), .RN(n3042), .Q(
        \CACHE[7][147] ), .QN(n1773) );
  DFFRX1 \CACHE_reg[7][146]  ( .D(n3012), .CK(clk), .RN(n3043), .Q(
        \CACHE[7][146] ), .QN(n1772) );
  DFFRX1 \CACHE_reg[7][145]  ( .D(n3011), .CK(clk), .RN(n3044), .Q(
        \CACHE[7][145] ), .QN(n1771) );
  DFFRX1 \CACHE_reg[7][144]  ( .D(n3010), .CK(clk), .RN(n3044), .Q(
        \CACHE[7][144] ), .QN(n1770) );
  DFFRX1 \CACHE_reg[7][143]  ( .D(n3009), .CK(clk), .RN(n3045), .Q(
        \CACHE[7][143] ), .QN(n1769) );
  DFFRX1 \CACHE_reg[7][142]  ( .D(n3008), .CK(clk), .RN(n3046), .Q(
        \CACHE[7][142] ), .QN(n1768) );
  DFFRX1 \CACHE_reg[7][141]  ( .D(n3007), .CK(clk), .RN(n3046), .Q(
        \CACHE[7][141] ), .QN(n1767) );
  DFFRX1 \CACHE_reg[7][140]  ( .D(n3006), .CK(clk), .RN(n3047), .Q(
        \CACHE[7][140] ), .QN(n1766) );
  DFFRX1 \CACHE_reg[7][139]  ( .D(n3005), .CK(clk), .RN(n3048), .Q(
        \CACHE[7][139] ), .QN(n1765) );
  DFFRX1 \CACHE_reg[7][138]  ( .D(n3004), .CK(clk), .RN(n3048), .Q(
        \CACHE[7][138] ), .QN(n1764) );
  DFFRX1 \CACHE_reg[7][137]  ( .D(n3003), .CK(clk), .RN(n3049), .Q(
        \CACHE[7][137] ), .QN(n1763) );
  DFFRX1 \CACHE_reg[7][136]  ( .D(n3002), .CK(clk), .RN(n3050), .Q(
        \CACHE[7][136] ), .QN(n1762) );
  DFFRX1 \CACHE_reg[7][135]  ( .D(n3001), .CK(clk), .RN(n3050), .Q(
        \CACHE[7][135] ), .QN(n1761) );
  DFFRX1 \CACHE_reg[7][134]  ( .D(n3000), .CK(clk), .RN(n3051), .Q(
        \CACHE[7][134] ), .QN(n1760) );
  DFFRX1 \CACHE_reg[7][133]  ( .D(n2999), .CK(clk), .RN(n3052), .Q(
        \CACHE[7][133] ), .QN(n1759) );
  DFFRX1 \CACHE_reg[7][132]  ( .D(n2998), .CK(clk), .RN(n3052), .Q(
        \CACHE[7][132] ), .QN(n1758) );
  DFFRX1 \CACHE_reg[7][131]  ( .D(n2997), .CK(clk), .RN(n3053), .Q(
        \CACHE[7][131] ), .QN(n1757) );
  DFFRX1 \CACHE_reg[7][130]  ( .D(n2996), .CK(clk), .RN(n3054), .Q(
        \CACHE[7][130] ), .QN(n1756) );
  DFFRX1 \CACHE_reg[7][129]  ( .D(n2995), .CK(clk), .RN(n3054), .Q(
        \CACHE[7][129] ), .QN(n1755) );
  DFFRX1 \CACHE_reg[7][128]  ( .D(n2994), .CK(clk), .RN(n3055), .Q(
        \CACHE[7][128] ), .QN(n1754) );
  DFFRX1 \CACHE_reg[7][127]  ( .D(n2993), .CK(clk), .RN(n478), .Q(
        \CACHE[7][127] ), .QN(n1753) );
  DFFRX1 \CACHE_reg[7][126]  ( .D(n2992), .CK(clk), .RN(n480), .Q(
        \CACHE[7][126] ), .QN(n1752) );
  DFFRX1 \CACHE_reg[7][125]  ( .D(n2991), .CK(clk), .RN(n483), .Q(
        \CACHE[7][125] ), .QN(n1751) );
  DFFRX1 \CACHE_reg[7][124]  ( .D(n2990), .CK(clk), .RN(n486), .Q(
        \CACHE[7][124] ), .QN(n1750) );
  DFFRX1 \CACHE_reg[7][123]  ( .D(n2989), .CK(clk), .RN(n488), .Q(
        \CACHE[7][123] ), .QN(n1749) );
  DFFRX1 \CACHE_reg[7][122]  ( .D(n2988), .CK(clk), .RN(n491), .Q(
        \CACHE[7][122] ), .QN(n1748) );
  DFFRX1 \CACHE_reg[7][121]  ( .D(n2987), .CK(clk), .RN(n494), .Q(
        \CACHE[7][121] ), .QN(n1747) );
  DFFRX1 \CACHE_reg[7][120]  ( .D(n2986), .CK(clk), .RN(n496), .Q(
        \CACHE[7][120] ), .QN(n1746) );
  DFFRX1 \CACHE_reg[7][119]  ( .D(n2985), .CK(clk), .RN(n499), .Q(
        \CACHE[7][119] ), .QN(n1745) );
  DFFRX1 \CACHE_reg[7][118]  ( .D(n2984), .CK(clk), .RN(n502), .Q(
        \CACHE[7][118] ), .QN(n1744) );
  DFFRX1 \CACHE_reg[7][117]  ( .D(n2983), .CK(clk), .RN(n504), .Q(
        \CACHE[7][117] ), .QN(n1743) );
  DFFRX1 \CACHE_reg[7][116]  ( .D(n2982), .CK(clk), .RN(n507), .Q(
        \CACHE[7][116] ), .QN(n1742) );
  DFFRX1 \CACHE_reg[7][115]  ( .D(n2981), .CK(clk), .RN(n510), .Q(
        \CACHE[7][115] ), .QN(n1741) );
  DFFRX1 \CACHE_reg[7][114]  ( .D(n2980), .CK(clk), .RN(n3033), .Q(
        \CACHE[7][114] ), .QN(n1740) );
  DFFRX1 \CACHE_reg[7][113]  ( .D(n2979), .CK(clk), .RN(n512), .Q(
        \CACHE[7][113] ), .QN(n1739) );
  DFFRX1 \CACHE_reg[7][112]  ( .D(n2978), .CK(clk), .RN(n515), .Q(
        \CACHE[7][112] ), .QN(n1738) );
  DFFRX1 \CACHE_reg[7][111]  ( .D(n2977), .CK(clk), .RN(n518), .Q(
        \CACHE[7][111] ), .QN(n1737) );
  DFFRX1 \CACHE_reg[7][110]  ( .D(n2976), .CK(clk), .RN(n520), .Q(
        \CACHE[7][110] ), .QN(n1736) );
  DFFRX1 \CACHE_reg[7][109]  ( .D(n2975), .CK(clk), .RN(n523), .Q(
        \CACHE[7][109] ), .QN(n1735) );
  DFFRX1 \CACHE_reg[7][108]  ( .D(n2974), .CK(clk), .RN(n526), .Q(
        \CACHE[7][108] ), .QN(n1734) );
  DFFRX1 \CACHE_reg[7][107]  ( .D(n2973), .CK(clk), .RN(n528), .Q(
        \CACHE[7][107] ), .QN(n1733) );
  DFFRX1 \CACHE_reg[7][106]  ( .D(n2972), .CK(clk), .RN(n531), .Q(
        \CACHE[7][106] ), .QN(n1732) );
  DFFRX1 \CACHE_reg[7][105]  ( .D(n2971), .CK(clk), .RN(n534), .Q(
        \CACHE[7][105] ), .QN(n1731) );
  DFFRX1 \CACHE_reg[7][104]  ( .D(n2970), .CK(clk), .RN(n536), .Q(
        \CACHE[7][104] ), .QN(n1730) );
  DFFRX1 \CACHE_reg[7][103]  ( .D(n2969), .CK(clk), .RN(n539), .Q(
        \CACHE[7][103] ), .QN(n1729) );
  DFFRX1 \CACHE_reg[7][102]  ( .D(n2968), .CK(clk), .RN(n3022), .Q(
        \CACHE[7][102] ), .QN(n1728) );
  DFFRX1 \CACHE_reg[7][101]  ( .D(n2967), .CK(clk), .RN(n3024), .Q(
        \CACHE[7][101] ), .QN(n1727) );
  DFFRX1 \CACHE_reg[7][100]  ( .D(n2966), .CK(clk), .RN(n3034), .Q(
        \CACHE[7][100] ), .QN(n1726) );
  DFFRX1 \CACHE_reg[7][99]  ( .D(n2965), .CK(clk), .RN(n3027), .Q(
        \CACHE[7][99] ), .QN(n1725) );
  DFFRX1 \CACHE_reg[7][98]  ( .D(n2964), .CK(clk), .RN(n3030), .Q(
        \CACHE[7][98] ), .QN(n1724) );
  DFFRX1 \CACHE_reg[7][97]  ( .D(n2963), .CK(clk), .RN(n3034), .Q(
        \CACHE[7][97] ), .QN(n1723) );
  DFFRX1 \CACHE_reg[7][96]  ( .D(n2962), .CK(clk), .RN(n3032), .Q(
        \CACHE[7][96] ), .QN(n1722) );
  DFFRX1 \CACHE_reg[7][95]  ( .D(n2961), .CK(clk), .RN(n477), .Q(
        \CACHE[7][95] ), .QN(n1721) );
  DFFRX1 \CACHE_reg[7][94]  ( .D(n2960), .CK(clk), .RN(n480), .Q(
        \CACHE[7][94] ), .QN(n1720) );
  DFFRX1 \CACHE_reg[7][93]  ( .D(n2959), .CK(clk), .RN(n482), .Q(
        \CACHE[7][93] ), .QN(n1719) );
  DFFRX1 \CACHE_reg[7][92]  ( .D(n2958), .CK(clk), .RN(n485), .Q(
        \CACHE[7][92] ), .QN(n1718) );
  DFFRX1 \CACHE_reg[7][91]  ( .D(n2957), .CK(clk), .RN(n488), .Q(
        \CACHE[7][91] ), .QN(n1717) );
  DFFRX1 \CACHE_reg[7][90]  ( .D(n2956), .CK(clk), .RN(n490), .Q(
        \CACHE[7][90] ), .QN(n1716) );
  DFFRX1 \CACHE_reg[7][89]  ( .D(n2955), .CK(clk), .RN(n493), .Q(
        \CACHE[7][89] ), .QN(n1715) );
  DFFRX1 \CACHE_reg[7][88]  ( .D(n2954), .CK(clk), .RN(n496), .Q(
        \CACHE[7][88] ), .QN(n1714) );
  DFFRX1 \CACHE_reg[7][87]  ( .D(n2953), .CK(clk), .RN(n498), .Q(
        \CACHE[7][87] ), .QN(n1713) );
  DFFRX1 \CACHE_reg[7][86]  ( .D(n2952), .CK(clk), .RN(n501), .Q(
        \CACHE[7][86] ), .QN(n1712) );
  DFFRX1 \CACHE_reg[7][85]  ( .D(n2951), .CK(clk), .RN(n504), .Q(
        \CACHE[7][85] ), .QN(n1711) );
  DFFRX1 \CACHE_reg[7][84]  ( .D(n2950), .CK(clk), .RN(n506), .Q(
        \CACHE[7][84] ), .QN(n1710) );
  DFFRX1 \CACHE_reg[7][83]  ( .D(n2949), .CK(clk), .RN(n509), .Q(
        \CACHE[7][83] ), .QN(n1709) );
  DFFRX1 \CACHE_reg[7][82]  ( .D(n2948), .CK(clk), .RN(n3035), .Q(
        \CACHE[7][82] ), .QN(n1708) );
  DFFRX1 \CACHE_reg[7][81]  ( .D(n2947), .CK(clk), .RN(n512), .Q(
        \CACHE[7][81] ), .QN(n1707) );
  DFFRX1 \CACHE_reg[7][80]  ( .D(n2946), .CK(clk), .RN(n514), .Q(
        \CACHE[7][80] ), .QN(n1706) );
  DFFRX1 \CACHE_reg[7][79]  ( .D(n2945), .CK(clk), .RN(n517), .Q(
        \CACHE[7][79] ), .QN(n1705) );
  DFFRX1 \CACHE_reg[7][78]  ( .D(n2944), .CK(clk), .RN(n520), .Q(
        \CACHE[7][78] ), .QN(n1704) );
  DFFRX1 \CACHE_reg[7][77]  ( .D(n2943), .CK(clk), .RN(n522), .Q(
        \CACHE[7][77] ), .QN(n1703) );
  DFFRX1 \CACHE_reg[7][76]  ( .D(n2942), .CK(clk), .RN(n525), .Q(
        \CACHE[7][76] ), .QN(n1702) );
  DFFRX1 \CACHE_reg[7][75]  ( .D(n2941), .CK(clk), .RN(n528), .Q(
        \CACHE[7][75] ), .QN(n1701) );
  DFFRX1 \CACHE_reg[7][74]  ( .D(n2940), .CK(clk), .RN(n530), .Q(
        \CACHE[7][74] ), .QN(n1700) );
  DFFRX1 \CACHE_reg[7][73]  ( .D(n2939), .CK(clk), .RN(n533), .Q(
        \CACHE[7][73] ), .QN(n1699) );
  DFFRX1 \CACHE_reg[7][72]  ( .D(n2938), .CK(clk), .RN(n536), .Q(
        \CACHE[7][72] ), .QN(n1698) );
  DFFRX1 \CACHE_reg[7][71]  ( .D(n2937), .CK(clk), .RN(n538), .Q(
        \CACHE[7][71] ), .QN(n1697) );
  DFFRX1 \CACHE_reg[7][70]  ( .D(n2936), .CK(clk), .RN(n3020), .Q(
        \CACHE[7][70] ), .QN(n1696) );
  DFFRX1 \CACHE_reg[7][69]  ( .D(n2935), .CK(clk), .RN(n3024), .Q(
        \CACHE[7][69] ), .QN(n1695) );
  DFFRX1 \CACHE_reg[7][68]  ( .D(n2934), .CK(clk), .RN(n3036), .Q(
        \CACHE[7][68] ), .QN(n1694) );
  DFFRX1 \CACHE_reg[7][67]  ( .D(n2933), .CK(clk), .RN(n3026), .Q(
        \CACHE[7][67] ), .QN(n1693) );
  DFFRX1 \CACHE_reg[7][66]  ( .D(n2932), .CK(clk), .RN(n3029), .Q(
        \CACHE[7][66] ), .QN(n1692) );
  DFFRX1 \CACHE_reg[7][65]  ( .D(n2931), .CK(clk), .RN(n3036), .Q(
        \CACHE[7][65] ), .QN(n1691) );
  DFFRX1 \CACHE_reg[7][64]  ( .D(n2930), .CK(clk), .RN(n3032), .Q(
        \CACHE[7][64] ), .QN(n1690) );
  DFFRX1 \CACHE_reg[7][63]  ( .D(n2929), .CK(clk), .RN(n476), .Q(
        \CACHE[7][63] ), .QN(n1689) );
  DFFRX1 \CACHE_reg[7][62]  ( .D(n2928), .CK(clk), .RN(n479), .Q(
        \CACHE[7][62] ), .QN(n1688) );
  DFFRX1 \CACHE_reg[7][61]  ( .D(n2927), .CK(clk), .RN(n482), .Q(
        \CACHE[7][61] ), .QN(n1687) );
  DFFRX1 \CACHE_reg[7][60]  ( .D(n2926), .CK(clk), .RN(n484), .Q(
        \CACHE[7][60] ), .QN(n1686) );
  DFFRX1 \CACHE_reg[7][59]  ( .D(n2925), .CK(clk), .RN(n487), .Q(
        \CACHE[7][59] ), .QN(n1685) );
  DFFRX1 \CACHE_reg[7][58]  ( .D(n2924), .CK(clk), .RN(n490), .Q(
        \CACHE[7][58] ), .QN(n1684) );
  DFFRX1 \CACHE_reg[7][57]  ( .D(n2923), .CK(clk), .RN(n492), .Q(
        \CACHE[7][57] ), .QN(n1683) );
  DFFRX1 \CACHE_reg[7][56]  ( .D(n2922), .CK(clk), .RN(n495), .Q(
        \CACHE[7][56] ), .QN(n1682) );
  DFFRX1 \CACHE_reg[7][55]  ( .D(n2921), .CK(clk), .RN(n498), .Q(
        \CACHE[7][55] ), .QN(n1681) );
  DFFRX1 \CACHE_reg[7][54]  ( .D(n2920), .CK(clk), .RN(n500), .Q(
        \CACHE[7][54] ), .QN(n1680) );
  DFFRX1 \CACHE_reg[7][53]  ( .D(n2919), .CK(clk), .RN(n503), .Q(
        \CACHE[7][53] ), .QN(n1679) );
  DFFRX1 \CACHE_reg[7][52]  ( .D(n2918), .CK(clk), .RN(n506), .Q(
        \CACHE[7][52] ), .QN(n1678) );
  DFFRX1 \CACHE_reg[7][51]  ( .D(n2917), .CK(clk), .RN(n508), .Q(
        \CACHE[7][51] ), .QN(n1677) );
  DFFRX1 \CACHE_reg[7][50]  ( .D(n2916), .CK(clk), .RN(n3037), .Q(
        \CACHE[7][50] ), .QN(n1676) );
  DFFRX1 \CACHE_reg[7][49]  ( .D(n2915), .CK(clk), .RN(n511), .Q(
        \CACHE[7][49] ), .QN(n1675) );
  DFFRX1 \CACHE_reg[7][48]  ( .D(n2914), .CK(clk), .RN(n514), .Q(
        \CACHE[7][48] ), .QN(n1674) );
  DFFRX1 \CACHE_reg[7][47]  ( .D(n2913), .CK(clk), .RN(n516), .Q(
        \CACHE[7][47] ), .QN(n1673) );
  DFFRX1 \CACHE_reg[7][46]  ( .D(n2912), .CK(clk), .RN(n519), .Q(
        \CACHE[7][46] ), .QN(n1672) );
  DFFRX1 \CACHE_reg[7][45]  ( .D(n2911), .CK(clk), .RN(n522), .Q(
        \CACHE[7][45] ), .QN(n1671) );
  DFFRX1 \CACHE_reg[7][44]  ( .D(n2910), .CK(clk), .RN(n524), .Q(
        \CACHE[7][44] ), .QN(n1670) );
  DFFRX1 \CACHE_reg[7][43]  ( .D(n2909), .CK(clk), .RN(n527), .Q(
        \CACHE[7][43] ), .QN(n1669) );
  DFFRX1 \CACHE_reg[7][42]  ( .D(n2908), .CK(clk), .RN(n530), .Q(
        \CACHE[7][42] ), .QN(n1668) );
  DFFRX1 \CACHE_reg[7][41]  ( .D(n2907), .CK(clk), .RN(n532), .Q(
        \CACHE[7][41] ), .QN(n1667) );
  DFFRX1 \CACHE_reg[7][40]  ( .D(n2906), .CK(clk), .RN(n535), .Q(
        \CACHE[7][40] ), .QN(n1666) );
  DFFRX1 \CACHE_reg[7][39]  ( .D(n2905), .CK(clk), .RN(n538), .Q(
        \CACHE[7][39] ), .QN(n1665) );
  DFFRX1 \CACHE_reg[7][38]  ( .D(n2904), .CK(clk), .RN(n540), .Q(
        \CACHE[7][38] ), .QN(n1664) );
  DFFRX1 \CACHE_reg[7][37]  ( .D(n2903), .CK(clk), .RN(n3023), .Q(
        \CACHE[7][37] ), .QN(n1663) );
  DFFRX1 \CACHE_reg[7][36]  ( .D(n2902), .CK(clk), .RN(n3038), .Q(
        \CACHE[7][36] ), .QN(n1662) );
  DFFRX1 \CACHE_reg[7][35]  ( .D(n2901), .CK(clk), .RN(n3026), .Q(
        \CACHE[7][35] ), .QN(n1661) );
  DFFRX1 \CACHE_reg[7][34]  ( .D(n2900), .CK(clk), .RN(n3028), .Q(
        \CACHE[7][34] ), .QN(n1660) );
  DFFRX1 \CACHE_reg[7][33]  ( .D(n2899), .CK(clk), .RN(n3038), .Q(
        \CACHE[7][33] ), .QN(n1659) );
  DFFRX1 \CACHE_reg[7][32]  ( .D(n2898), .CK(clk), .RN(n3031), .Q(
        \CACHE[7][32] ), .QN(n1658) );
  DFFRX1 \CACHE_reg[7][31]  ( .D(n2897), .CK(clk), .RN(n476), .Q(
        \CACHE[7][31] ), .QN(n1657) );
  DFFRX1 \CACHE_reg[7][30]  ( .D(n2896), .CK(clk), .RN(n478), .Q(
        \CACHE[7][30] ), .QN(n1656) );
  DFFRX1 \CACHE_reg[7][29]  ( .D(n2895), .CK(clk), .RN(n481), .Q(
        \CACHE[7][29] ), .QN(n1655) );
  DFFRX1 \CACHE_reg[7][28]  ( .D(n2894), .CK(clk), .RN(n484), .Q(
        \CACHE[7][28] ), .QN(n1654) );
  DFFRX1 \CACHE_reg[7][27]  ( .D(n2893), .CK(clk), .RN(n486), .Q(
        \CACHE[7][27] ), .QN(n1653) );
  DFFRX1 \CACHE_reg[7][26]  ( .D(n2892), .CK(clk), .RN(n489), .Q(
        \CACHE[7][26] ), .QN(n1652) );
  DFFRX1 \CACHE_reg[7][25]  ( .D(n2891), .CK(clk), .RN(n492), .Q(
        \CACHE[7][25] ), .QN(n1651) );
  DFFRX1 \CACHE_reg[7][24]  ( .D(n2890), .CK(clk), .RN(n494), .Q(
        \CACHE[7][24] ), .QN(n1650) );
  DFFRX1 \CACHE_reg[7][23]  ( .D(n2889), .CK(clk), .RN(n497), .Q(
        \CACHE[7][23] ), .QN(n1649) );
  DFFRX1 \CACHE_reg[7][22]  ( .D(n2888), .CK(clk), .RN(n500), .Q(
        \CACHE[7][22] ), .QN(n1648) );
  DFFRX1 \CACHE_reg[7][21]  ( .D(n2887), .CK(clk), .RN(n502), .Q(
        \CACHE[7][21] ), .QN(n1647) );
  DFFRX1 \CACHE_reg[7][20]  ( .D(n2886), .CK(clk), .RN(n505), .Q(
        \CACHE[7][20] ), .QN(n1646) );
  DFFRX1 \CACHE_reg[7][19]  ( .D(n2885), .CK(clk), .RN(n508), .Q(
        \CACHE[7][19] ), .QN(n1645) );
  DFFRX1 \CACHE_reg[7][18]  ( .D(n2884), .CK(clk), .RN(n3058), .Q(
        \CACHE[7][18] ), .QN(n1644) );
  DFFRX1 \CACHE_reg[7][17]  ( .D(n2883), .CK(clk), .RN(n510), .Q(
        \CACHE[7][17] ), .QN(n1643) );
  DFFRX1 \CACHE_reg[7][16]  ( .D(n2882), .CK(clk), .RN(n513), .Q(
        \CACHE[7][16] ), .QN(n1642) );
  DFFRX1 \CACHE_reg[7][15]  ( .D(n2881), .CK(clk), .RN(n516), .Q(
        \CACHE[7][15] ), .QN(n1641) );
  DFFRX1 \CACHE_reg[7][14]  ( .D(n2880), .CK(clk), .RN(n518), .Q(
        \CACHE[7][14] ), .QN(n1640) );
  DFFRX1 \CACHE_reg[7][13]  ( .D(n2879), .CK(clk), .RN(n521), .Q(
        \CACHE[7][13] ), .QN(n1639) );
  DFFRX1 \CACHE_reg[7][12]  ( .D(n2878), .CK(clk), .RN(n524), .Q(
        \CACHE[7][12] ), .QN(n1638) );
  DFFRX1 \CACHE_reg[7][11]  ( .D(n2877), .CK(clk), .RN(n526), .Q(
        \CACHE[7][11] ), .QN(n1637) );
  DFFRX1 \CACHE_reg[7][10]  ( .D(n2876), .CK(clk), .RN(n529), .Q(
        \CACHE[7][10] ), .QN(n1636) );
  DFFRX1 \CACHE_reg[7][9]  ( .D(n2875), .CK(clk), .RN(n532), .Q(\CACHE[7][9] ), 
        .QN(n1635) );
  DFFRX1 \CACHE_reg[7][8]  ( .D(n2874), .CK(clk), .RN(n534), .Q(\CACHE[7][8] ), 
        .QN(n1634) );
  DFFRX1 \CACHE_reg[7][7]  ( .D(n2873), .CK(clk), .RN(n537), .Q(\CACHE[7][7] ), 
        .QN(n1633) );
  DFFRX1 \CACHE_reg[7][6]  ( .D(n2872), .CK(clk), .RN(n540), .Q(\CACHE[7][6] ), 
        .QN(n1632) );
  DFFRX1 \CACHE_reg[7][5]  ( .D(n2871), .CK(clk), .RN(n3022), .Q(\CACHE[7][5] ), .QN(n1631) );
  DFFRX1 \CACHE_reg[7][4]  ( .D(n2870), .CK(clk), .RN(n3058), .Q(\CACHE[7][4] ), .QN(n1630) );
  DFFRX1 \CACHE_reg[7][3]  ( .D(n2869), .CK(clk), .RN(n3025), .Q(\CACHE[7][3] ), .QN(n1629) );
  DFFRX1 \CACHE_reg[7][2]  ( .D(n2868), .CK(clk), .RN(n3028), .Q(\CACHE[7][2] ), .QN(n1628) );
  DFFRX1 \CACHE_reg[7][1]  ( .D(n2867), .CK(clk), .RN(n3039), .Q(\CACHE[7][1] ), .QN(n1627) );
  DFFRX1 \CACHE_reg[7][0]  ( .D(n2866), .CK(clk), .RN(n3030), .Q(\CACHE[7][0] ), .QN(n1626) );
  DFFRX1 \CACHE_reg[3][154]  ( .D(n2400), .CK(clk), .RN(n3057), .Q(
        \CACHE[3][154] ), .QN(n1160) );
  DFFRX1 \CACHE_reg[3][153]  ( .D(n2399), .CK(clk), .RN(n3057), .Q(
        \CACHE[3][153] ), .QN(n1159) );
  DFFRX1 \CACHE_reg[3][152]  ( .D(n2398), .CK(clk), .RN(n3056), .Q(
        \CACHE[3][152] ), .QN(n1158) );
  DFFRX1 \CACHE_reg[3][151]  ( .D(n2397), .CK(clk), .RN(n3040), .Q(
        \CACHE[3][151] ), .QN(n1157) );
  DFFRX1 \CACHE_reg[3][150]  ( .D(n2396), .CK(clk), .RN(n3041), .Q(
        \CACHE[3][150] ), .QN(n1156) );
  DFFRX1 \CACHE_reg[3][149]  ( .D(n2395), .CK(clk), .RN(n3041), .Q(
        \CACHE[3][149] ), .QN(n1155) );
  DFFRX1 \CACHE_reg[3][148]  ( .D(n2394), .CK(clk), .RN(n3042), .Q(
        \CACHE[3][148] ), .QN(n1154) );
  DFFRX1 \CACHE_reg[3][147]  ( .D(n2393), .CK(clk), .RN(n3043), .Q(
        \CACHE[3][147] ), .QN(n1153) );
  DFFRX1 \CACHE_reg[3][146]  ( .D(n2392), .CK(clk), .RN(n3043), .Q(
        \CACHE[3][146] ), .QN(n1152) );
  DFFRX1 \CACHE_reg[3][145]  ( .D(n2391), .CK(clk), .RN(n3044), .Q(
        \CACHE[3][145] ), .QN(n1151) );
  DFFRX1 \CACHE_reg[3][144]  ( .D(n2390), .CK(clk), .RN(n3045), .Q(
        \CACHE[3][144] ), .QN(n1150) );
  DFFRX1 \CACHE_reg[3][143]  ( .D(n2389), .CK(clk), .RN(n3045), .Q(
        \CACHE[3][143] ), .QN(n1149) );
  DFFRX1 \CACHE_reg[3][142]  ( .D(n2388), .CK(clk), .RN(n3046), .Q(
        \CACHE[3][142] ), .QN(n1148) );
  DFFRX1 \CACHE_reg[3][141]  ( .D(n2387), .CK(clk), .RN(n3047), .Q(
        \CACHE[3][141] ), .QN(n1147) );
  DFFRX1 \CACHE_reg[3][140]  ( .D(n2386), .CK(clk), .RN(n3047), .Q(
        \CACHE[3][140] ), .QN(n1146) );
  DFFRX1 \CACHE_reg[3][139]  ( .D(n2385), .CK(clk), .RN(n3048), .Q(
        \CACHE[3][139] ), .QN(n1145) );
  DFFRX1 \CACHE_reg[3][138]  ( .D(n2384), .CK(clk), .RN(n3049), .Q(
        \CACHE[3][138] ), .QN(n1144) );
  DFFRX1 \CACHE_reg[3][137]  ( .D(n2383), .CK(clk), .RN(n3049), .Q(
        \CACHE[3][137] ), .QN(n1143) );
  DFFRX1 \CACHE_reg[3][136]  ( .D(n2382), .CK(clk), .RN(n3050), .Q(
        \CACHE[3][136] ), .QN(n1142) );
  DFFRX1 \CACHE_reg[3][135]  ( .D(n2381), .CK(clk), .RN(n3051), .Q(
        \CACHE[3][135] ), .QN(n1141) );
  DFFRX1 \CACHE_reg[3][134]  ( .D(n2380), .CK(clk), .RN(n3051), .Q(
        \CACHE[3][134] ), .QN(n1140) );
  DFFRX1 \CACHE_reg[3][133]  ( .D(n2379), .CK(clk), .RN(n3052), .Q(
        \CACHE[3][133] ), .QN(n1139) );
  DFFRX1 \CACHE_reg[3][132]  ( .D(n2378), .CK(clk), .RN(n3053), .Q(
        \CACHE[3][132] ), .QN(n1138) );
  DFFRX1 \CACHE_reg[3][131]  ( .D(n2377), .CK(clk), .RN(n3053), .Q(
        \CACHE[3][131] ), .QN(n1137) );
  DFFRX1 \CACHE_reg[3][130]  ( .D(n2376), .CK(clk), .RN(n3054), .Q(
        \CACHE[3][130] ), .QN(n1136) );
  DFFRX1 \CACHE_reg[3][129]  ( .D(n2375), .CK(clk), .RN(n3055), .Q(
        \CACHE[3][129] ), .QN(n1135) );
  DFFRX1 \CACHE_reg[3][128]  ( .D(n2374), .CK(clk), .RN(n3055), .Q(
        \CACHE[3][128] ), .QN(n1134) );
  DFFRX1 \CACHE_reg[3][127]  ( .D(n2373), .CK(clk), .RN(n478), .Q(
        \CACHE[3][127] ), .QN(n1133) );
  DFFRX1 \CACHE_reg[3][126]  ( .D(n2372), .CK(clk), .RN(n481), .Q(
        \CACHE[3][126] ), .QN(n1132) );
  DFFRX1 \CACHE_reg[3][125]  ( .D(n2371), .CK(clk), .RN(n483), .Q(
        \CACHE[3][125] ), .QN(n1131) );
  DFFRX1 \CACHE_reg[3][124]  ( .D(n2370), .CK(clk), .RN(n486), .Q(
        \CACHE[3][124] ), .QN(n1130) );
  DFFRX1 \CACHE_reg[3][123]  ( .D(n2369), .CK(clk), .RN(n489), .Q(
        \CACHE[3][123] ), .QN(n1129) );
  DFFRX1 \CACHE_reg[3][122]  ( .D(n2368), .CK(clk), .RN(n491), .Q(
        \CACHE[3][122] ), .QN(n1128) );
  DFFRX1 \CACHE_reg[3][121]  ( .D(n2367), .CK(clk), .RN(n494), .Q(
        \CACHE[3][121] ), .QN(n1127) );
  DFFRX1 \CACHE_reg[3][120]  ( .D(n2366), .CK(clk), .RN(n497), .Q(
        \CACHE[3][120] ), .QN(n1126) );
  DFFRX1 \CACHE_reg[3][119]  ( .D(n2365), .CK(clk), .RN(n499), .Q(
        \CACHE[3][119] ), .QN(n1125) );
  DFFRX1 \CACHE_reg[3][118]  ( .D(n2364), .CK(clk), .RN(n502), .Q(
        \CACHE[3][118] ), .QN(n1124) );
  DFFRX1 \CACHE_reg[3][117]  ( .D(n2363), .CK(clk), .RN(n505), .Q(
        \CACHE[3][117] ), .QN(n1123) );
  DFFRX1 \CACHE_reg[3][116]  ( .D(n2362), .CK(clk), .RN(n507), .Q(
        \CACHE[3][116] ), .QN(n1122) );
  DFFRX1 \CACHE_reg[3][115]  ( .D(n2361), .CK(clk), .RN(n510), .Q(
        \CACHE[3][115] ), .QN(n1121) );
  DFFRX1 \CACHE_reg[3][114]  ( .D(n2360), .CK(clk), .RN(n3033), .Q(
        \CACHE[3][114] ), .QN(n1120) );
  DFFRX1 \CACHE_reg[3][113]  ( .D(n2359), .CK(clk), .RN(n513), .Q(
        \CACHE[3][113] ), .QN(n1119) );
  DFFRX1 \CACHE_reg[3][112]  ( .D(n2358), .CK(clk), .RN(n515), .Q(
        \CACHE[3][112] ), .QN(n1118) );
  DFFRX1 \CACHE_reg[3][111]  ( .D(n2357), .CK(clk), .RN(n518), .Q(
        \CACHE[3][111] ), .QN(n1117) );
  DFFRX1 \CACHE_reg[3][110]  ( .D(n2356), .CK(clk), .RN(n521), .Q(
        \CACHE[3][110] ), .QN(n1116) );
  DFFRX1 \CACHE_reg[3][109]  ( .D(n2355), .CK(clk), .RN(n523), .Q(
        \CACHE[3][109] ), .QN(n1115) );
  DFFRX1 \CACHE_reg[3][108]  ( .D(n2354), .CK(clk), .RN(n526), .Q(
        \CACHE[3][108] ), .QN(n1114) );
  DFFRX1 \CACHE_reg[3][107]  ( .D(n2353), .CK(clk), .RN(n529), .Q(
        \CACHE[3][107] ), .QN(n1113) );
  DFFRX1 \CACHE_reg[3][106]  ( .D(n2352), .CK(clk), .RN(n531), .Q(
        \CACHE[3][106] ), .QN(n1112) );
  DFFRX1 \CACHE_reg[3][105]  ( .D(n2351), .CK(clk), .RN(n534), .Q(
        \CACHE[3][105] ), .QN(n1111) );
  DFFRX1 \CACHE_reg[3][104]  ( .D(n2350), .CK(clk), .RN(n537), .Q(
        \CACHE[3][104] ), .QN(n1110) );
  DFFRX1 \CACHE_reg[3][103]  ( .D(n2349), .CK(clk), .RN(n539), .Q(
        \CACHE[3][103] ), .QN(n1109) );
  DFFRX1 \CACHE_reg[3][102]  ( .D(n2348), .CK(clk), .RN(n3022), .Q(
        \CACHE[3][102] ), .QN(n1108) );
  DFFRX1 \CACHE_reg[3][101]  ( .D(n2347), .CK(clk), .RN(n3025), .Q(
        \CACHE[3][101] ), .QN(n1107) );
  DFFRX1 \CACHE_reg[3][100]  ( .D(n2346), .CK(clk), .RN(n3034), .Q(
        \CACHE[3][100] ), .QN(n1106) );
  DFFRX1 \CACHE_reg[3][99]  ( .D(n2345), .CK(clk), .RN(n3027), .Q(
        \CACHE[3][99] ), .QN(n1105) );
  DFFRX1 \CACHE_reg[3][98]  ( .D(n2344), .CK(clk), .RN(n3030), .Q(
        \CACHE[3][98] ), .QN(n1104) );
  DFFRX1 \CACHE_reg[3][97]  ( .D(n2343), .CK(clk), .RN(n3035), .Q(
        \CACHE[3][97] ), .QN(n1103) );
  DFFRX1 \CACHE_reg[3][96]  ( .D(n2342), .CK(clk), .RN(n3033), .Q(
        \CACHE[3][96] ), .QN(n1102) );
  DFFRX1 \CACHE_reg[3][95]  ( .D(n2341), .CK(clk), .RN(n477), .Q(
        \CACHE[3][95] ), .QN(n1101) );
  DFFRX1 \CACHE_reg[3][94]  ( .D(n2340), .CK(clk), .RN(n480), .Q(
        \CACHE[3][94] ), .QN(n1100) );
  DFFRX1 \CACHE_reg[3][93]  ( .D(n2339), .CK(clk), .RN(n483), .Q(
        \CACHE[3][93] ), .QN(n1099) );
  DFFRX1 \CACHE_reg[3][92]  ( .D(n2338), .CK(clk), .RN(n485), .Q(
        \CACHE[3][92] ), .QN(n1098) );
  DFFRX1 \CACHE_reg[3][91]  ( .D(n2337), .CK(clk), .RN(n488), .Q(
        \CACHE[3][91] ), .QN(n1097) );
  DFFRX1 \CACHE_reg[3][90]  ( .D(n2336), .CK(clk), .RN(n491), .Q(
        \CACHE[3][90] ), .QN(n1096) );
  DFFRX1 \CACHE_reg[3][89]  ( .D(n2335), .CK(clk), .RN(n493), .Q(
        \CACHE[3][89] ), .QN(n1095) );
  DFFRX1 \CACHE_reg[3][88]  ( .D(n2334), .CK(clk), .RN(n496), .Q(
        \CACHE[3][88] ), .QN(n1094) );
  DFFRX1 \CACHE_reg[3][87]  ( .D(n2333), .CK(clk), .RN(n499), .Q(
        \CACHE[3][87] ), .QN(n1093) );
  DFFRX1 \CACHE_reg[3][86]  ( .D(n2332), .CK(clk), .RN(n501), .Q(
        \CACHE[3][86] ), .QN(n1092) );
  DFFRX1 \CACHE_reg[3][85]  ( .D(n2331), .CK(clk), .RN(n504), .Q(
        \CACHE[3][85] ), .QN(n1091) );
  DFFRX1 \CACHE_reg[3][84]  ( .D(n2330), .CK(clk), .RN(n507), .Q(
        \CACHE[3][84] ), .QN(n1090) );
  DFFRX1 \CACHE_reg[3][83]  ( .D(n2329), .CK(clk), .RN(n509), .Q(
        \CACHE[3][83] ), .QN(n1089) );
  DFFRX1 \CACHE_reg[3][82]  ( .D(n2328), .CK(clk), .RN(n3035), .Q(
        \CACHE[3][82] ), .QN(n1088) );
  DFFRX1 \CACHE_reg[3][81]  ( .D(n2327), .CK(clk), .RN(n512), .Q(
        \CACHE[3][81] ), .QN(n1087) );
  DFFRX1 \CACHE_reg[3][80]  ( .D(n2326), .CK(clk), .RN(n515), .Q(
        \CACHE[3][80] ), .QN(n1086) );
  DFFRX1 \CACHE_reg[3][79]  ( .D(n2325), .CK(clk), .RN(n517), .Q(
        \CACHE[3][79] ), .QN(n1085) );
  DFFRX1 \CACHE_reg[3][78]  ( .D(n2324), .CK(clk), .RN(n520), .Q(
        \CACHE[3][78] ), .QN(n1084) );
  DFFRX1 \CACHE_reg[3][77]  ( .D(n2323), .CK(clk), .RN(n523), .Q(
        \CACHE[3][77] ), .QN(n1083) );
  DFFRX1 \CACHE_reg[3][76]  ( .D(n2322), .CK(clk), .RN(n525), .Q(
        \CACHE[3][76] ), .QN(n1082) );
  DFFRX1 \CACHE_reg[3][75]  ( .D(n2321), .CK(clk), .RN(n528), .Q(
        \CACHE[3][75] ), .QN(n1081) );
  DFFRX1 \CACHE_reg[3][74]  ( .D(n2320), .CK(clk), .RN(n531), .Q(
        \CACHE[3][74] ), .QN(n1080) );
  DFFRX1 \CACHE_reg[3][73]  ( .D(n2319), .CK(clk), .RN(n533), .Q(
        \CACHE[3][73] ), .QN(n1079) );
  DFFRX1 \CACHE_reg[3][72]  ( .D(n2318), .CK(clk), .RN(n536), .Q(
        \CACHE[3][72] ), .QN(n1078) );
  DFFRX1 \CACHE_reg[3][71]  ( .D(n2317), .CK(clk), .RN(n539), .Q(
        \CACHE[3][71] ), .QN(n1077) );
  DFFRX1 \CACHE_reg[3][70]  ( .D(n2316), .CK(clk), .RN(n3020), .Q(
        \CACHE[3][70] ), .QN(n1076) );
  DFFRX1 \CACHE_reg[3][69]  ( .D(n2315), .CK(clk), .RN(n3024), .Q(
        \CACHE[3][69] ), .QN(n1075) );
  DFFRX1 \CACHE_reg[3][68]  ( .D(n2314), .CK(clk), .RN(n3036), .Q(
        \CACHE[3][68] ), .QN(n1074) );
  DFFRX1 \CACHE_reg[3][67]  ( .D(n2313), .CK(clk), .RN(n3027), .Q(
        \CACHE[3][67] ), .QN(n1073) );
  DFFRX1 \CACHE_reg[3][66]  ( .D(n2312), .CK(clk), .RN(n3029), .Q(
        \CACHE[3][66] ), .QN(n1072) );
  DFFRX1 \CACHE_reg[3][65]  ( .D(n2311), .CK(clk), .RN(n3037), .Q(
        \CACHE[3][65] ), .QN(n1071) );
  DFFRX1 \CACHE_reg[3][64]  ( .D(n2310), .CK(clk), .RN(n3032), .Q(
        \CACHE[3][64] ), .QN(n1070) );
  DFFRX1 \CACHE_reg[3][63]  ( .D(n2309), .CK(clk), .RN(n477), .Q(
        \CACHE[3][63] ), .QN(n1069) );
  DFFRX1 \CACHE_reg[3][62]  ( .D(n2308), .CK(clk), .RN(n479), .Q(
        \CACHE[3][62] ), .QN(n1068) );
  DFFRX1 \CACHE_reg[3][61]  ( .D(n2307), .CK(clk), .RN(n482), .Q(
        \CACHE[3][61] ), .QN(n1067) );
  DFFRX1 \CACHE_reg[3][60]  ( .D(n2306), .CK(clk), .RN(n485), .Q(
        \CACHE[3][60] ), .QN(n1066) );
  DFFRX1 \CACHE_reg[3][59]  ( .D(n2305), .CK(clk), .RN(n487), .Q(
        \CACHE[3][59] ), .QN(n1065) );
  DFFRX1 \CACHE_reg[3][58]  ( .D(n2304), .CK(clk), .RN(n490), .Q(
        \CACHE[3][58] ), .QN(n1064) );
  DFFRX1 \CACHE_reg[3][57]  ( .D(n2303), .CK(clk), .RN(n493), .Q(
        \CACHE[3][57] ), .QN(n1063) );
  DFFRX1 \CACHE_reg[3][56]  ( .D(n2302), .CK(clk), .RN(n495), .Q(
        \CACHE[3][56] ), .QN(n1062) );
  DFFRX1 \CACHE_reg[3][55]  ( .D(n2301), .CK(clk), .RN(n498), .Q(
        \CACHE[3][55] ), .QN(n1061) );
  DFFRX1 \CACHE_reg[3][54]  ( .D(n2300), .CK(clk), .RN(n501), .Q(
        \CACHE[3][54] ), .QN(n1060) );
  DFFRX1 \CACHE_reg[3][53]  ( .D(n2299), .CK(clk), .RN(n503), .Q(
        \CACHE[3][53] ), .QN(n1059) );
  DFFRX1 \CACHE_reg[3][52]  ( .D(n2298), .CK(clk), .RN(n506), .Q(
        \CACHE[3][52] ), .QN(n1058) );
  DFFRX1 \CACHE_reg[3][51]  ( .D(n2297), .CK(clk), .RN(n509), .Q(
        \CACHE[3][51] ), .QN(n1057) );
  DFFRX1 \CACHE_reg[3][50]  ( .D(n2296), .CK(clk), .RN(n3037), .Q(
        \CACHE[3][50] ), .QN(n1056) );
  DFFRX1 \CACHE_reg[3][49]  ( .D(n2295), .CK(clk), .RN(n511), .Q(
        \CACHE[3][49] ), .QN(n1055) );
  DFFRX1 \CACHE_reg[3][48]  ( .D(n2294), .CK(clk), .RN(n514), .Q(
        \CACHE[3][48] ), .QN(n1054) );
  DFFRX1 \CACHE_reg[3][47]  ( .D(n2293), .CK(clk), .RN(n517), .Q(
        \CACHE[3][47] ), .QN(n1053) );
  DFFRX1 \CACHE_reg[3][46]  ( .D(n2292), .CK(clk), .RN(n519), .Q(
        \CACHE[3][46] ), .QN(n1052) );
  DFFRX1 \CACHE_reg[3][45]  ( .D(n2291), .CK(clk), .RN(n522), .Q(
        \CACHE[3][45] ), .QN(n1051) );
  DFFRX1 \CACHE_reg[3][44]  ( .D(n2290), .CK(clk), .RN(n525), .Q(
        \CACHE[3][44] ), .QN(n1050) );
  DFFRX1 \CACHE_reg[3][43]  ( .D(n2289), .CK(clk), .RN(n527), .Q(
        \CACHE[3][43] ), .QN(n1049) );
  DFFRX1 \CACHE_reg[3][42]  ( .D(n2288), .CK(clk), .RN(n530), .Q(
        \CACHE[3][42] ), .QN(n1048) );
  DFFRX1 \CACHE_reg[3][41]  ( .D(n2287), .CK(clk), .RN(n533), .Q(
        \CACHE[3][41] ), .QN(n1047) );
  DFFRX1 \CACHE_reg[3][40]  ( .D(n2286), .CK(clk), .RN(n535), .Q(
        \CACHE[3][40] ), .QN(n1046) );
  DFFRX1 \CACHE_reg[3][39]  ( .D(n2285), .CK(clk), .RN(n538), .Q(
        \CACHE[3][39] ), .QN(n1045) );
  DFFRX1 \CACHE_reg[3][38]  ( .D(n2284), .CK(clk), .RN(n3020), .Q(
        \CACHE[3][38] ), .QN(n1044) );
  DFFRX1 \CACHE_reg[3][37]  ( .D(n2283), .CK(clk), .RN(n3023), .Q(
        \CACHE[3][37] ), .QN(n1043) );
  DFFRX1 \CACHE_reg[3][36]  ( .D(n2282), .CK(clk), .RN(n3038), .Q(
        \CACHE[3][36] ), .QN(n1042) );
  DFFRX1 \CACHE_reg[3][35]  ( .D(n2281), .CK(clk), .RN(n3026), .Q(
        \CACHE[3][35] ), .QN(n1041) );
  DFFRX1 \CACHE_reg[3][34]  ( .D(n2280), .CK(clk), .RN(n3029), .Q(
        \CACHE[3][34] ), .QN(n1040) );
  DFFRX1 \CACHE_reg[3][33]  ( .D(n2279), .CK(clk), .RN(n3039), .Q(
        \CACHE[3][33] ), .QN(n1039) );
  DFFRX1 \CACHE_reg[3][32]  ( .D(n2278), .CK(clk), .RN(n3031), .Q(
        \CACHE[3][32] ), .QN(n1038) );
  DFFRX1 \CACHE_reg[3][31]  ( .D(n2277), .CK(clk), .RN(n476), .Q(
        \CACHE[3][31] ), .QN(n1037) );
  DFFRX1 \CACHE_reg[3][30]  ( .D(n2276), .CK(clk), .RN(n479), .Q(
        \CACHE[3][30] ), .QN(n1036) );
  DFFRX1 \CACHE_reg[3][29]  ( .D(n2275), .CK(clk), .RN(n481), .Q(
        \CACHE[3][29] ), .QN(n1035) );
  DFFRX1 \CACHE_reg[3][28]  ( .D(n2274), .CK(clk), .RN(n484), .Q(
        \CACHE[3][28] ), .QN(n1034) );
  DFFRX1 \CACHE_reg[3][27]  ( .D(n2273), .CK(clk), .RN(n487), .Q(
        \CACHE[3][27] ), .QN(n1033) );
  DFFRX1 \CACHE_reg[3][26]  ( .D(n2272), .CK(clk), .RN(n489), .Q(
        \CACHE[3][26] ), .QN(n1032) );
  DFFRX1 \CACHE_reg[3][25]  ( .D(n2271), .CK(clk), .RN(n492), .Q(
        \CACHE[3][25] ), .QN(n1031) );
  DFFRX1 \CACHE_reg[3][24]  ( .D(n2270), .CK(clk), .RN(n495), .Q(
        \CACHE[3][24] ), .QN(n1030) );
  DFFRX1 \CACHE_reg[3][23]  ( .D(n2269), .CK(clk), .RN(n497), .Q(
        \CACHE[3][23] ), .QN(n1029) );
  DFFRX1 \CACHE_reg[3][22]  ( .D(n2268), .CK(clk), .RN(n500), .Q(
        \CACHE[3][22] ), .QN(n1028) );
  DFFRX1 \CACHE_reg[3][21]  ( .D(n2267), .CK(clk), .RN(n503), .Q(
        \CACHE[3][21] ), .QN(n1027) );
  DFFRX1 \CACHE_reg[3][20]  ( .D(n2266), .CK(clk), .RN(n505), .Q(
        \CACHE[3][20] ), .QN(n1026) );
  DFFRX1 \CACHE_reg[3][19]  ( .D(n2265), .CK(clk), .RN(n508), .Q(
        \CACHE[3][19] ), .QN(n1025) );
  DFFRX1 \CACHE_reg[3][18]  ( .D(n2264), .CK(clk), .RN(n3059), .Q(
        \CACHE[3][18] ), .QN(n1024) );
  DFFRX1 \CACHE_reg[3][17]  ( .D(n2263), .CK(clk), .RN(n511), .Q(
        \CACHE[3][17] ), .QN(n1023) );
  DFFRX1 \CACHE_reg[3][16]  ( .D(n2262), .CK(clk), .RN(n513), .Q(
        \CACHE[3][16] ), .QN(n1022) );
  DFFRX1 \CACHE_reg[3][15]  ( .D(n2261), .CK(clk), .RN(n516), .Q(
        \CACHE[3][15] ), .QN(n1021) );
  DFFRX1 \CACHE_reg[3][14]  ( .D(n2260), .CK(clk), .RN(n519), .Q(
        \CACHE[3][14] ), .QN(n1020) );
  DFFRX1 \CACHE_reg[3][13]  ( .D(n2259), .CK(clk), .RN(n521), .Q(
        \CACHE[3][13] ), .QN(n1019) );
  DFFRX1 \CACHE_reg[3][12]  ( .D(n2258), .CK(clk), .RN(n524), .Q(
        \CACHE[3][12] ), .QN(n1018) );
  DFFRX1 \CACHE_reg[3][11]  ( .D(n2257), .CK(clk), .RN(n527), .Q(
        \CACHE[3][11] ), .QN(n1017) );
  DFFRX1 \CACHE_reg[3][10]  ( .D(n2256), .CK(clk), .RN(n529), .Q(
        \CACHE[3][10] ), .QN(n1016) );
  DFFRX1 \CACHE_reg[3][9]  ( .D(n2255), .CK(clk), .RN(n532), .Q(\CACHE[3][9] ), 
        .QN(n1015) );
  DFFRX1 \CACHE_reg[3][8]  ( .D(n2254), .CK(clk), .RN(n535), .Q(\CACHE[3][8] ), 
        .QN(n1014) );
  DFFRX1 \CACHE_reg[3][7]  ( .D(n2253), .CK(clk), .RN(n537), .Q(\CACHE[3][7] ), 
        .QN(n1013) );
  DFFRX1 \CACHE_reg[3][6]  ( .D(n2252), .CK(clk), .RN(n540), .Q(\CACHE[3][6] ), 
        .QN(n1012) );
  DFFRX1 \CACHE_reg[3][5]  ( .D(n2251), .CK(clk), .RN(n3023), .Q(\CACHE[3][5] ), .QN(n1011) );
  DFFRX1 \CACHE_reg[3][4]  ( .D(n2250), .CK(clk), .RN(n3058), .Q(\CACHE[3][4] ), .QN(n1010) );
  DFFRX1 \CACHE_reg[3][3]  ( .D(n2249), .CK(clk), .RN(n3025), .Q(\CACHE[3][3] ), .QN(n1009) );
  DFFRX1 \CACHE_reg[3][2]  ( .D(n2248), .CK(clk), .RN(n3028), .Q(\CACHE[3][2] ), .QN(n1008) );
  DFFRX1 \CACHE_reg[3][1]  ( .D(n2247), .CK(clk), .RN(n3039), .Q(\CACHE[3][1] ), .QN(n1007) );
  DFFRX1 \CACHE_reg[3][0]  ( .D(n2246), .CK(clk), .RN(n3031), .Q(\CACHE[3][0] ), .QN(n1006) );
  DFFRX1 \CACHE_reg[5][154]  ( .D(n2710), .CK(clk), .RN(n3057), .Q(
        \CACHE[5][154] ), .QN(n1470) );
  DFFRX1 \CACHE_reg[5][153]  ( .D(n2709), .CK(clk), .RN(n3056), .Q(
        \CACHE[5][153] ), .QN(n1469) );
  DFFRX1 \CACHE_reg[5][152]  ( .D(n2708), .CK(clk), .RN(n3056), .Q(
        \CACHE[5][152] ), .QN(n1468) );
  DFFRX1 \CACHE_reg[5][151]  ( .D(n2707), .CK(clk), .RN(n3040), .Q(
        \CACHE[5][151] ), .QN(n1467) );
  DFFRX1 \CACHE_reg[5][150]  ( .D(n2706), .CK(clk), .RN(n3040), .Q(
        \CACHE[5][150] ), .QN(n1466) );
  DFFRX1 \CACHE_reg[5][149]  ( .D(n2705), .CK(clk), .RN(n3041), .Q(
        \CACHE[5][149] ), .QN(n1465) );
  DFFRX1 \CACHE_reg[5][148]  ( .D(n2704), .CK(clk), .RN(n3042), .Q(
        \CACHE[5][148] ), .QN(n1464) );
  DFFRX1 \CACHE_reg[5][147]  ( .D(n2703), .CK(clk), .RN(n3042), .Q(
        \CACHE[5][147] ), .QN(n1463) );
  DFFRX1 \CACHE_reg[5][146]  ( .D(n2702), .CK(clk), .RN(n3043), .Q(
        \CACHE[5][146] ), .QN(n1462) );
  DFFRX1 \CACHE_reg[5][145]  ( .D(n2701), .CK(clk), .RN(n3044), .Q(
        \CACHE[5][145] ), .QN(n1461) );
  DFFRX1 \CACHE_reg[5][144]  ( .D(n2700), .CK(clk), .RN(n3044), .Q(
        \CACHE[5][144] ), .QN(n1460) );
  DFFRX1 \CACHE_reg[5][143]  ( .D(n2699), .CK(clk), .RN(n3045), .Q(
        \CACHE[5][143] ), .QN(n1459) );
  DFFRX1 \CACHE_reg[5][142]  ( .D(n2698), .CK(clk), .RN(n3046), .Q(
        \CACHE[5][142] ), .QN(n1458) );
  DFFRX1 \CACHE_reg[5][141]  ( .D(n2697), .CK(clk), .RN(n3046), .Q(
        \CACHE[5][141] ), .QN(n1457) );
  DFFRX1 \CACHE_reg[5][140]  ( .D(n2696), .CK(clk), .RN(n3047), .Q(
        \CACHE[5][140] ), .QN(n1456) );
  DFFRX1 \CACHE_reg[5][139]  ( .D(n2695), .CK(clk), .RN(n3048), .Q(
        \CACHE[5][139] ), .QN(n1455) );
  DFFRX1 \CACHE_reg[5][138]  ( .D(n2694), .CK(clk), .RN(n3048), .Q(
        \CACHE[5][138] ), .QN(n1454) );
  DFFRX1 \CACHE_reg[5][137]  ( .D(n2693), .CK(clk), .RN(n3049), .Q(
        \CACHE[5][137] ), .QN(n1453) );
  DFFRX1 \CACHE_reg[5][136]  ( .D(n2692), .CK(clk), .RN(n3050), .Q(
        \CACHE[5][136] ), .QN(n1452) );
  DFFRX1 \CACHE_reg[5][135]  ( .D(n2691), .CK(clk), .RN(n3050), .Q(
        \CACHE[5][135] ), .QN(n1451) );
  DFFRX1 \CACHE_reg[5][134]  ( .D(n2690), .CK(clk), .RN(n3051), .Q(
        \CACHE[5][134] ), .QN(n1450) );
  DFFRX1 \CACHE_reg[5][133]  ( .D(n2689), .CK(clk), .RN(n3052), .Q(
        \CACHE[5][133] ), .QN(n1449) );
  DFFRX1 \CACHE_reg[5][132]  ( .D(n2688), .CK(clk), .RN(n3052), .Q(
        \CACHE[5][132] ), .QN(n1448) );
  DFFRX1 \CACHE_reg[5][131]  ( .D(n2687), .CK(clk), .RN(n3053), .Q(
        \CACHE[5][131] ), .QN(n1447) );
  DFFRX1 \CACHE_reg[5][130]  ( .D(n2686), .CK(clk), .RN(n3054), .Q(
        \CACHE[5][130] ), .QN(n1446) );
  DFFRX1 \CACHE_reg[5][129]  ( .D(n2685), .CK(clk), .RN(n3054), .Q(
        \CACHE[5][129] ), .QN(n1445) );
  DFFRX1 \CACHE_reg[5][128]  ( .D(n2684), .CK(clk), .RN(n3055), .Q(
        \CACHE[5][128] ), .QN(n1444) );
  DFFRX1 \CACHE_reg[5][127]  ( .D(n2683), .CK(clk), .RN(n478), .Q(
        \CACHE[5][127] ), .QN(n1443) );
  DFFRX1 \CACHE_reg[5][126]  ( .D(n2682), .CK(clk), .RN(n480), .Q(
        \CACHE[5][126] ), .QN(n1442) );
  DFFRX1 \CACHE_reg[5][125]  ( .D(n2681), .CK(clk), .RN(n483), .Q(
        \CACHE[5][125] ), .QN(n1441) );
  DFFRX1 \CACHE_reg[5][124]  ( .D(n2680), .CK(clk), .RN(n486), .Q(
        \CACHE[5][124] ), .QN(n1440) );
  DFFRX1 \CACHE_reg[5][123]  ( .D(n2679), .CK(clk), .RN(n488), .Q(
        \CACHE[5][123] ), .QN(n1439) );
  DFFRX1 \CACHE_reg[5][122]  ( .D(n2678), .CK(clk), .RN(n491), .Q(
        \CACHE[5][122] ), .QN(n1438) );
  DFFRX1 \CACHE_reg[5][121]  ( .D(n2677), .CK(clk), .RN(n494), .Q(
        \CACHE[5][121] ), .QN(n1437) );
  DFFRX1 \CACHE_reg[5][120]  ( .D(n2676), .CK(clk), .RN(n496), .Q(
        \CACHE[5][120] ), .QN(n1436) );
  DFFRX1 \CACHE_reg[5][119]  ( .D(n2675), .CK(clk), .RN(n499), .Q(
        \CACHE[5][119] ), .QN(n1435) );
  DFFRX1 \CACHE_reg[5][118]  ( .D(n2674), .CK(clk), .RN(n502), .Q(
        \CACHE[5][118] ), .QN(n1434) );
  DFFRX1 \CACHE_reg[5][117]  ( .D(n2673), .CK(clk), .RN(n504), .Q(
        \CACHE[5][117] ), .QN(n1433) );
  DFFRX1 \CACHE_reg[5][116]  ( .D(n2672), .CK(clk), .RN(n507), .Q(
        \CACHE[5][116] ), .QN(n1432) );
  DFFRX1 \CACHE_reg[5][115]  ( .D(n2671), .CK(clk), .RN(n510), .Q(
        \CACHE[5][115] ), .QN(n1431) );
  DFFRX1 \CACHE_reg[5][114]  ( .D(n2670), .CK(clk), .RN(n3033), .Q(
        \CACHE[5][114] ), .QN(n1430) );
  DFFRX1 \CACHE_reg[5][113]  ( .D(n2669), .CK(clk), .RN(n512), .Q(
        \CACHE[5][113] ), .QN(n1429) );
  DFFRX1 \CACHE_reg[5][112]  ( .D(n2668), .CK(clk), .RN(n515), .Q(
        \CACHE[5][112] ), .QN(n1428) );
  DFFRX1 \CACHE_reg[5][111]  ( .D(n2667), .CK(clk), .RN(n518), .Q(
        \CACHE[5][111] ), .QN(n1427) );
  DFFRX1 \CACHE_reg[5][110]  ( .D(n2666), .CK(clk), .RN(n520), .Q(
        \CACHE[5][110] ), .QN(n1426) );
  DFFRX1 \CACHE_reg[5][109]  ( .D(n2665), .CK(clk), .RN(n523), .Q(
        \CACHE[5][109] ), .QN(n1425) );
  DFFRX1 \CACHE_reg[5][108]  ( .D(n2664), .CK(clk), .RN(n526), .Q(
        \CACHE[5][108] ), .QN(n1424) );
  DFFRX1 \CACHE_reg[5][107]  ( .D(n2663), .CK(clk), .RN(n528), .Q(
        \CACHE[5][107] ), .QN(n1423) );
  DFFRX1 \CACHE_reg[5][106]  ( .D(n2662), .CK(clk), .RN(n531), .Q(
        \CACHE[5][106] ), .QN(n1422) );
  DFFRX1 \CACHE_reg[5][105]  ( .D(n2661), .CK(clk), .RN(n534), .Q(
        \CACHE[5][105] ), .QN(n1421) );
  DFFRX1 \CACHE_reg[5][104]  ( .D(n2660), .CK(clk), .RN(n536), .Q(
        \CACHE[5][104] ), .QN(n1420) );
  DFFRX1 \CACHE_reg[5][103]  ( .D(n2659), .CK(clk), .RN(n539), .Q(
        \CACHE[5][103] ), .QN(n1419) );
  DFFRX1 \CACHE_reg[5][102]  ( .D(n2658), .CK(clk), .RN(n3022), .Q(
        \CACHE[5][102] ), .QN(n1418) );
  DFFRX1 \CACHE_reg[5][101]  ( .D(n2657), .CK(clk), .RN(n3024), .Q(
        \CACHE[5][101] ), .QN(n1417) );
  DFFRX1 \CACHE_reg[5][100]  ( .D(n2656), .CK(clk), .RN(n3034), .Q(
        \CACHE[5][100] ), .QN(n1416) );
  DFFRX1 \CACHE_reg[5][99]  ( .D(n2655), .CK(clk), .RN(n3027), .Q(
        \CACHE[5][99] ), .QN(n1415) );
  DFFRX1 \CACHE_reg[5][98]  ( .D(n2654), .CK(clk), .RN(n3030), .Q(
        \CACHE[5][98] ), .QN(n1414) );
  DFFRX1 \CACHE_reg[5][97]  ( .D(n2653), .CK(clk), .RN(n3034), .Q(
        \CACHE[5][97] ), .QN(n1413) );
  DFFRX1 \CACHE_reg[5][96]  ( .D(n2652), .CK(clk), .RN(n3032), .Q(
        \CACHE[5][96] ), .QN(n1412) );
  DFFRX1 \CACHE_reg[5][95]  ( .D(n2651), .CK(clk), .RN(n477), .Q(
        \CACHE[5][95] ), .QN(n1411) );
  DFFRX1 \CACHE_reg[5][94]  ( .D(n2650), .CK(clk), .RN(n480), .Q(
        \CACHE[5][94] ), .QN(n1410) );
  DFFRX1 \CACHE_reg[5][93]  ( .D(n2649), .CK(clk), .RN(n482), .Q(
        \CACHE[5][93] ), .QN(n1409) );
  DFFRX1 \CACHE_reg[5][92]  ( .D(n2648), .CK(clk), .RN(n485), .Q(
        \CACHE[5][92] ), .QN(n1408) );
  DFFRX1 \CACHE_reg[5][91]  ( .D(n2647), .CK(clk), .RN(n488), .Q(
        \CACHE[5][91] ), .QN(n1407) );
  DFFRX1 \CACHE_reg[5][90]  ( .D(n2646), .CK(clk), .RN(n490), .Q(
        \CACHE[5][90] ), .QN(n1406) );
  DFFRX1 \CACHE_reg[5][89]  ( .D(n2645), .CK(clk), .RN(n493), .Q(
        \CACHE[5][89] ), .QN(n1405) );
  DFFRX1 \CACHE_reg[5][88]  ( .D(n2644), .CK(clk), .RN(n496), .Q(
        \CACHE[5][88] ), .QN(n1404) );
  DFFRX1 \CACHE_reg[5][87]  ( .D(n2643), .CK(clk), .RN(n498), .Q(
        \CACHE[5][87] ), .QN(n1403) );
  DFFRX1 \CACHE_reg[5][86]  ( .D(n2642), .CK(clk), .RN(n501), .Q(
        \CACHE[5][86] ), .QN(n1402) );
  DFFRX1 \CACHE_reg[5][85]  ( .D(n2641), .CK(clk), .RN(n504), .Q(
        \CACHE[5][85] ), .QN(n1401) );
  DFFRX1 \CACHE_reg[5][84]  ( .D(n2640), .CK(clk), .RN(n506), .Q(
        \CACHE[5][84] ), .QN(n1400) );
  DFFRX1 \CACHE_reg[5][83]  ( .D(n2639), .CK(clk), .RN(n509), .Q(
        \CACHE[5][83] ), .QN(n1399) );
  DFFRX1 \CACHE_reg[5][82]  ( .D(n2638), .CK(clk), .RN(n3035), .Q(
        \CACHE[5][82] ), .QN(n1398) );
  DFFRX1 \CACHE_reg[5][81]  ( .D(n2637), .CK(clk), .RN(n512), .Q(
        \CACHE[5][81] ), .QN(n1397) );
  DFFRX1 \CACHE_reg[5][80]  ( .D(n2636), .CK(clk), .RN(n514), .Q(
        \CACHE[5][80] ), .QN(n1396) );
  DFFRX1 \CACHE_reg[5][79]  ( .D(n2635), .CK(clk), .RN(n517), .Q(
        \CACHE[5][79] ), .QN(n1395) );
  DFFRX1 \CACHE_reg[5][78]  ( .D(n2634), .CK(clk), .RN(n520), .Q(
        \CACHE[5][78] ), .QN(n1394) );
  DFFRX1 \CACHE_reg[5][77]  ( .D(n2633), .CK(clk), .RN(n522), .Q(
        \CACHE[5][77] ), .QN(n1393) );
  DFFRX1 \CACHE_reg[5][76]  ( .D(n2632), .CK(clk), .RN(n525), .Q(
        \CACHE[5][76] ), .QN(n1392) );
  DFFRX1 \CACHE_reg[5][75]  ( .D(n2631), .CK(clk), .RN(n528), .Q(
        \CACHE[5][75] ), .QN(n1391) );
  DFFRX1 \CACHE_reg[5][74]  ( .D(n2630), .CK(clk), .RN(n530), .Q(
        \CACHE[5][74] ), .QN(n1390) );
  DFFRX1 \CACHE_reg[5][73]  ( .D(n2629), .CK(clk), .RN(n533), .Q(
        \CACHE[5][73] ), .QN(n1389) );
  DFFRX1 \CACHE_reg[5][72]  ( .D(n2628), .CK(clk), .RN(n536), .Q(
        \CACHE[5][72] ), .QN(n1388) );
  DFFRX1 \CACHE_reg[5][71]  ( .D(n2627), .CK(clk), .RN(n538), .Q(
        \CACHE[5][71] ), .QN(n1387) );
  DFFRX1 \CACHE_reg[5][70]  ( .D(n2626), .CK(clk), .RN(n3020), .Q(
        \CACHE[5][70] ), .QN(n1386) );
  DFFRX1 \CACHE_reg[5][69]  ( .D(n2625), .CK(clk), .RN(n3024), .Q(
        \CACHE[5][69] ), .QN(n1385) );
  DFFRX1 \CACHE_reg[5][68]  ( .D(n2624), .CK(clk), .RN(n3036), .Q(
        \CACHE[5][68] ), .QN(n1384) );
  DFFRX1 \CACHE_reg[5][67]  ( .D(n2623), .CK(clk), .RN(n3026), .Q(
        \CACHE[5][67] ), .QN(n1383) );
  DFFRX1 \CACHE_reg[5][66]  ( .D(n2622), .CK(clk), .RN(n3029), .Q(
        \CACHE[5][66] ), .QN(n1382) );
  DFFRX1 \CACHE_reg[5][65]  ( .D(n2621), .CK(clk), .RN(n3036), .Q(
        \CACHE[5][65] ), .QN(n1381) );
  DFFRX1 \CACHE_reg[5][64]  ( .D(n2620), .CK(clk), .RN(n3032), .Q(
        \CACHE[5][64] ), .QN(n1380) );
  DFFRX1 \CACHE_reg[5][63]  ( .D(n2619), .CK(clk), .RN(n476), .Q(
        \CACHE[5][63] ), .QN(n1379) );
  DFFRX1 \CACHE_reg[5][62]  ( .D(n2618), .CK(clk), .RN(n479), .Q(
        \CACHE[5][62] ), .QN(n1378) );
  DFFRX1 \CACHE_reg[5][61]  ( .D(n2617), .CK(clk), .RN(n482), .Q(
        \CACHE[5][61] ), .QN(n1377) );
  DFFRX1 \CACHE_reg[5][60]  ( .D(n2616), .CK(clk), .RN(n484), .Q(
        \CACHE[5][60] ), .QN(n1376) );
  DFFRX1 \CACHE_reg[5][59]  ( .D(n2615), .CK(clk), .RN(n487), .Q(
        \CACHE[5][59] ), .QN(n1375) );
  DFFRX1 \CACHE_reg[5][58]  ( .D(n2614), .CK(clk), .RN(n490), .Q(
        \CACHE[5][58] ), .QN(n1374) );
  DFFRX1 \CACHE_reg[5][57]  ( .D(n2613), .CK(clk), .RN(n492), .Q(
        \CACHE[5][57] ), .QN(n1373) );
  DFFRX1 \CACHE_reg[5][56]  ( .D(n2612), .CK(clk), .RN(n495), .Q(
        \CACHE[5][56] ), .QN(n1372) );
  DFFRX1 \CACHE_reg[5][55]  ( .D(n2611), .CK(clk), .RN(n498), .Q(
        \CACHE[5][55] ), .QN(n1371) );
  DFFRX1 \CACHE_reg[5][54]  ( .D(n2610), .CK(clk), .RN(n500), .Q(
        \CACHE[5][54] ), .QN(n1370) );
  DFFRX1 \CACHE_reg[5][53]  ( .D(n2609), .CK(clk), .RN(n503), .Q(
        \CACHE[5][53] ), .QN(n1369) );
  DFFRX1 \CACHE_reg[5][52]  ( .D(n2608), .CK(clk), .RN(n506), .Q(
        \CACHE[5][52] ), .QN(n1368) );
  DFFRX1 \CACHE_reg[5][51]  ( .D(n2607), .CK(clk), .RN(n508), .Q(
        \CACHE[5][51] ), .QN(n1367) );
  DFFRX1 \CACHE_reg[5][50]  ( .D(n2606), .CK(clk), .RN(n3037), .Q(
        \CACHE[5][50] ), .QN(n1366) );
  DFFRX1 \CACHE_reg[5][49]  ( .D(n2605), .CK(clk), .RN(n511), .Q(
        \CACHE[5][49] ), .QN(n1365) );
  DFFRX1 \CACHE_reg[5][48]  ( .D(n2604), .CK(clk), .RN(n514), .Q(
        \CACHE[5][48] ), .QN(n1364) );
  DFFRX1 \CACHE_reg[5][47]  ( .D(n2603), .CK(clk), .RN(n516), .Q(
        \CACHE[5][47] ), .QN(n1363) );
  DFFRX1 \CACHE_reg[5][46]  ( .D(n2602), .CK(clk), .RN(n519), .Q(
        \CACHE[5][46] ), .QN(n1362) );
  DFFRX1 \CACHE_reg[5][45]  ( .D(n2601), .CK(clk), .RN(n522), .Q(
        \CACHE[5][45] ), .QN(n1361) );
  DFFRX1 \CACHE_reg[5][44]  ( .D(n2600), .CK(clk), .RN(n524), .Q(
        \CACHE[5][44] ), .QN(n1360) );
  DFFRX1 \CACHE_reg[5][43]  ( .D(n2599), .CK(clk), .RN(n527), .Q(
        \CACHE[5][43] ), .QN(n1359) );
  DFFRX1 \CACHE_reg[5][42]  ( .D(n2598), .CK(clk), .RN(n530), .Q(
        \CACHE[5][42] ), .QN(n1358) );
  DFFRX1 \CACHE_reg[5][41]  ( .D(n2597), .CK(clk), .RN(n532), .Q(
        \CACHE[5][41] ), .QN(n1357) );
  DFFRX1 \CACHE_reg[5][40]  ( .D(n2596), .CK(clk), .RN(n535), .Q(
        \CACHE[5][40] ), .QN(n1356) );
  DFFRX1 \CACHE_reg[5][39]  ( .D(n2595), .CK(clk), .RN(n538), .Q(
        \CACHE[5][39] ), .QN(n1355) );
  DFFRX1 \CACHE_reg[5][38]  ( .D(n2594), .CK(clk), .RN(n540), .Q(
        \CACHE[5][38] ), .QN(n1354) );
  DFFRX1 \CACHE_reg[5][37]  ( .D(n2593), .CK(clk), .RN(n3023), .Q(
        \CACHE[5][37] ), .QN(n1353) );
  DFFRX1 \CACHE_reg[5][36]  ( .D(n2592), .CK(clk), .RN(n3038), .Q(
        \CACHE[5][36] ), .QN(n1352) );
  DFFRX1 \CACHE_reg[5][35]  ( .D(n2591), .CK(clk), .RN(n3026), .Q(
        \CACHE[5][35] ), .QN(n1351) );
  DFFRX1 \CACHE_reg[5][34]  ( .D(n2590), .CK(clk), .RN(n3028), .Q(
        \CACHE[5][34] ), .QN(n1350) );
  DFFRX1 \CACHE_reg[5][33]  ( .D(n2589), .CK(clk), .RN(n3038), .Q(
        \CACHE[5][33] ), .QN(n1349) );
  DFFRX1 \CACHE_reg[5][32]  ( .D(n2588), .CK(clk), .RN(n3031), .Q(
        \CACHE[5][32] ), .QN(n1348) );
  DFFRX1 \CACHE_reg[5][31]  ( .D(n2587), .CK(clk), .RN(n476), .Q(
        \CACHE[5][31] ), .QN(n1347) );
  DFFRX1 \CACHE_reg[5][30]  ( .D(n2586), .CK(clk), .RN(n478), .Q(
        \CACHE[5][30] ), .QN(n1346) );
  DFFRX1 \CACHE_reg[5][29]  ( .D(n2585), .CK(clk), .RN(n481), .Q(
        \CACHE[5][29] ), .QN(n1345) );
  DFFRX1 \CACHE_reg[5][28]  ( .D(n2584), .CK(clk), .RN(n484), .Q(
        \CACHE[5][28] ), .QN(n1344) );
  DFFRX1 \CACHE_reg[5][27]  ( .D(n2583), .CK(clk), .RN(n486), .Q(
        \CACHE[5][27] ), .QN(n1343) );
  DFFRX1 \CACHE_reg[5][26]  ( .D(n2582), .CK(clk), .RN(n489), .Q(
        \CACHE[5][26] ), .QN(n1342) );
  DFFRX1 \CACHE_reg[5][25]  ( .D(n2581), .CK(clk), .RN(n492), .Q(
        \CACHE[5][25] ), .QN(n1341) );
  DFFRX1 \CACHE_reg[5][24]  ( .D(n2580), .CK(clk), .RN(n494), .Q(
        \CACHE[5][24] ), .QN(n1340) );
  DFFRX1 \CACHE_reg[5][23]  ( .D(n2579), .CK(clk), .RN(n497), .Q(
        \CACHE[5][23] ), .QN(n1339) );
  DFFRX1 \CACHE_reg[5][22]  ( .D(n2578), .CK(clk), .RN(n500), .Q(
        \CACHE[5][22] ), .QN(n1338) );
  DFFRX1 \CACHE_reg[5][21]  ( .D(n2577), .CK(clk), .RN(n502), .Q(
        \CACHE[5][21] ), .QN(n1337) );
  DFFRX1 \CACHE_reg[5][20]  ( .D(n2576), .CK(clk), .RN(n505), .Q(
        \CACHE[5][20] ), .QN(n1336) );
  DFFRX1 \CACHE_reg[5][19]  ( .D(n2575), .CK(clk), .RN(n508), .Q(
        \CACHE[5][19] ), .QN(n1335) );
  DFFRX1 \CACHE_reg[5][18]  ( .D(n2574), .CK(clk), .RN(n3058), .Q(
        \CACHE[5][18] ), .QN(n1334) );
  DFFRX1 \CACHE_reg[5][17]  ( .D(n2573), .CK(clk), .RN(n510), .Q(
        \CACHE[5][17] ), .QN(n1333) );
  DFFRX1 \CACHE_reg[5][16]  ( .D(n2572), .CK(clk), .RN(n513), .Q(
        \CACHE[5][16] ), .QN(n1332) );
  DFFRX1 \CACHE_reg[5][15]  ( .D(n2571), .CK(clk), .RN(n516), .Q(
        \CACHE[5][15] ), .QN(n1331) );
  DFFRX1 \CACHE_reg[5][14]  ( .D(n2570), .CK(clk), .RN(n518), .Q(
        \CACHE[5][14] ), .QN(n1330) );
  DFFRX1 \CACHE_reg[5][13]  ( .D(n2569), .CK(clk), .RN(n521), .Q(
        \CACHE[5][13] ), .QN(n1329) );
  DFFRX1 \CACHE_reg[5][12]  ( .D(n2568), .CK(clk), .RN(n524), .Q(
        \CACHE[5][12] ), .QN(n1328) );
  DFFRX1 \CACHE_reg[5][11]  ( .D(n2567), .CK(clk), .RN(n526), .Q(
        \CACHE[5][11] ), .QN(n1327) );
  DFFRX1 \CACHE_reg[5][10]  ( .D(n2566), .CK(clk), .RN(n529), .Q(
        \CACHE[5][10] ), .QN(n1326) );
  DFFRX1 \CACHE_reg[5][9]  ( .D(n2565), .CK(clk), .RN(n532), .Q(\CACHE[5][9] ), 
        .QN(n1325) );
  DFFRX1 \CACHE_reg[5][8]  ( .D(n2564), .CK(clk), .RN(n534), .Q(\CACHE[5][8] ), 
        .QN(n1324) );
  DFFRX1 \CACHE_reg[5][7]  ( .D(n2563), .CK(clk), .RN(n537), .Q(\CACHE[5][7] ), 
        .QN(n1323) );
  DFFRX1 \CACHE_reg[5][6]  ( .D(n2562), .CK(clk), .RN(n540), .Q(\CACHE[5][6] ), 
        .QN(n1322) );
  DFFRX1 \CACHE_reg[5][5]  ( .D(n2561), .CK(clk), .RN(n3022), .Q(\CACHE[5][5] ), .QN(n1321) );
  DFFRX1 \CACHE_reg[5][4]  ( .D(n2560), .CK(clk), .RN(n3058), .Q(\CACHE[5][4] ), .QN(n1320) );
  DFFRX1 \CACHE_reg[5][3]  ( .D(n2559), .CK(clk), .RN(n3025), .Q(\CACHE[5][3] ), .QN(n1319) );
  DFFRX1 \CACHE_reg[5][2]  ( .D(n2558), .CK(clk), .RN(n3028), .Q(\CACHE[5][2] ), .QN(n1318) );
  DFFRX1 \CACHE_reg[5][1]  ( .D(n2557), .CK(clk), .RN(n3039), .Q(\CACHE[5][1] ), .QN(n1317) );
  DFFRX1 \CACHE_reg[5][0]  ( .D(n2556), .CK(clk), .RN(n3030), .Q(\CACHE[5][0] ), .QN(n1316) );
  DFFRX1 \CACHE_reg[1][154]  ( .D(n2090), .CK(clk), .RN(n3057), .Q(
        \CACHE[1][154] ), .QN(n850) );
  DFFRX1 \CACHE_reg[1][153]  ( .D(n2089), .CK(clk), .RN(n3057), .Q(
        \CACHE[1][153] ), .QN(n849) );
  DFFRX1 \CACHE_reg[1][152]  ( .D(n2088), .CK(clk), .RN(n3056), .Q(
        \CACHE[1][152] ), .QN(n848) );
  DFFRX1 \CACHE_reg[1][151]  ( .D(n2087), .CK(clk), .RN(n3040), .Q(
        \CACHE[1][151] ), .QN(n847) );
  DFFRX1 \CACHE_reg[1][150]  ( .D(n2086), .CK(clk), .RN(n3041), .Q(
        \CACHE[1][150] ), .QN(n846) );
  DFFRX1 \CACHE_reg[1][149]  ( .D(n2085), .CK(clk), .RN(n3041), .Q(
        \CACHE[1][149] ), .QN(n845) );
  DFFRX1 \CACHE_reg[1][148]  ( .D(n2084), .CK(clk), .RN(n3042), .Q(
        \CACHE[1][148] ), .QN(n844) );
  DFFRX1 \CACHE_reg[1][147]  ( .D(n2083), .CK(clk), .RN(n3043), .Q(
        \CACHE[1][147] ), .QN(n843) );
  DFFRX1 \CACHE_reg[1][146]  ( .D(n2082), .CK(clk), .RN(n3043), .Q(
        \CACHE[1][146] ), .QN(n842) );
  DFFRX1 \CACHE_reg[1][145]  ( .D(n2081), .CK(clk), .RN(n3044), .Q(
        \CACHE[1][145] ), .QN(n841) );
  DFFRX1 \CACHE_reg[1][144]  ( .D(n2080), .CK(clk), .RN(n3045), .Q(
        \CACHE[1][144] ), .QN(n840) );
  DFFRX1 \CACHE_reg[1][143]  ( .D(n2079), .CK(clk), .RN(n3045), .Q(
        \CACHE[1][143] ), .QN(n839) );
  DFFRX1 \CACHE_reg[1][142]  ( .D(n2078), .CK(clk), .RN(n3046), .Q(
        \CACHE[1][142] ), .QN(n838) );
  DFFRX1 \CACHE_reg[1][141]  ( .D(n2077), .CK(clk), .RN(n3047), .Q(
        \CACHE[1][141] ), .QN(n837) );
  DFFRX1 \CACHE_reg[1][140]  ( .D(n2076), .CK(clk), .RN(n3047), .Q(
        \CACHE[1][140] ), .QN(n836) );
  DFFRX1 \CACHE_reg[1][139]  ( .D(n2075), .CK(clk), .RN(n3048), .Q(
        \CACHE[1][139] ), .QN(n835) );
  DFFRX1 \CACHE_reg[1][138]  ( .D(n2074), .CK(clk), .RN(n3049), .Q(
        \CACHE[1][138] ), .QN(n834) );
  DFFRX1 \CACHE_reg[1][137]  ( .D(n2073), .CK(clk), .RN(n3049), .Q(
        \CACHE[1][137] ), .QN(n833) );
  DFFRX1 \CACHE_reg[1][136]  ( .D(n2072), .CK(clk), .RN(n3050), .Q(
        \CACHE[1][136] ), .QN(n832) );
  DFFRX1 \CACHE_reg[1][135]  ( .D(n2071), .CK(clk), .RN(n3051), .Q(
        \CACHE[1][135] ), .QN(n831) );
  DFFRX1 \CACHE_reg[1][134]  ( .D(n2070), .CK(clk), .RN(n3051), .Q(
        \CACHE[1][134] ), .QN(n830) );
  DFFRX1 \CACHE_reg[1][133]  ( .D(n2069), .CK(clk), .RN(n3052), .Q(
        \CACHE[1][133] ), .QN(n829) );
  DFFRX1 \CACHE_reg[1][132]  ( .D(n2068), .CK(clk), .RN(n3053), .Q(
        \CACHE[1][132] ), .QN(n828) );
  DFFRX1 \CACHE_reg[1][131]  ( .D(n2067), .CK(clk), .RN(n3053), .Q(
        \CACHE[1][131] ), .QN(n827) );
  DFFRX1 \CACHE_reg[1][130]  ( .D(n2066), .CK(clk), .RN(n3054), .Q(
        \CACHE[1][130] ), .QN(n826) );
  DFFRX1 \CACHE_reg[1][129]  ( .D(n2065), .CK(clk), .RN(n3055), .Q(
        \CACHE[1][129] ), .QN(n825) );
  DFFRX1 \CACHE_reg[1][128]  ( .D(n2064), .CK(clk), .RN(n3055), .Q(
        \CACHE[1][128] ), .QN(n824) );
  DFFRX1 \CACHE_reg[1][127]  ( .D(n2063), .CK(clk), .RN(n478), .Q(
        \CACHE[1][127] ), .QN(n823) );
  DFFRX1 \CACHE_reg[1][126]  ( .D(n2062), .CK(clk), .RN(n481), .Q(
        \CACHE[1][126] ), .QN(n822) );
  DFFRX1 \CACHE_reg[1][125]  ( .D(n2061), .CK(clk), .RN(n483), .Q(
        \CACHE[1][125] ), .QN(n821) );
  DFFRX1 \CACHE_reg[1][124]  ( .D(n2060), .CK(clk), .RN(n486), .Q(
        \CACHE[1][124] ), .QN(n820) );
  DFFRX1 \CACHE_reg[1][123]  ( .D(n2059), .CK(clk), .RN(n489), .Q(
        \CACHE[1][123] ), .QN(n819) );
  DFFRX1 \CACHE_reg[1][122]  ( .D(n2058), .CK(clk), .RN(n491), .Q(
        \CACHE[1][122] ), .QN(n818) );
  DFFRX1 \CACHE_reg[1][121]  ( .D(n2057), .CK(clk), .RN(n494), .Q(
        \CACHE[1][121] ), .QN(n817) );
  DFFRX1 \CACHE_reg[1][120]  ( .D(n2056), .CK(clk), .RN(n497), .Q(
        \CACHE[1][120] ), .QN(n816) );
  DFFRX1 \CACHE_reg[1][119]  ( .D(n2055), .CK(clk), .RN(n499), .Q(
        \CACHE[1][119] ), .QN(n815) );
  DFFRX1 \CACHE_reg[1][118]  ( .D(n2054), .CK(clk), .RN(n502), .Q(
        \CACHE[1][118] ), .QN(n814) );
  DFFRX1 \CACHE_reg[1][117]  ( .D(n2053), .CK(clk), .RN(n505), .Q(
        \CACHE[1][117] ), .QN(n813) );
  DFFRX1 \CACHE_reg[1][116]  ( .D(n2052), .CK(clk), .RN(n507), .Q(
        \CACHE[1][116] ), .QN(n812) );
  DFFRX1 \CACHE_reg[1][115]  ( .D(n2051), .CK(clk), .RN(n510), .Q(
        \CACHE[1][115] ), .QN(n811) );
  DFFRX1 \CACHE_reg[1][114]  ( .D(n2050), .CK(clk), .RN(n3033), .Q(
        \CACHE[1][114] ), .QN(n810) );
  DFFRX1 \CACHE_reg[1][113]  ( .D(n2049), .CK(clk), .RN(n513), .Q(
        \CACHE[1][113] ), .QN(n809) );
  DFFRX1 \CACHE_reg[1][112]  ( .D(n2048), .CK(clk), .RN(n515), .Q(
        \CACHE[1][112] ), .QN(n808) );
  DFFRX1 \CACHE_reg[1][111]  ( .D(n2047), .CK(clk), .RN(n518), .Q(
        \CACHE[1][111] ), .QN(n807) );
  DFFRX1 \CACHE_reg[1][110]  ( .D(n2046), .CK(clk), .RN(n521), .Q(
        \CACHE[1][110] ), .QN(n806) );
  DFFRX1 \CACHE_reg[1][109]  ( .D(n2045), .CK(clk), .RN(n523), .Q(
        \CACHE[1][109] ), .QN(n805) );
  DFFRX1 \CACHE_reg[1][108]  ( .D(n2044), .CK(clk), .RN(n526), .Q(
        \CACHE[1][108] ), .QN(n804) );
  DFFRX1 \CACHE_reg[1][107]  ( .D(n2043), .CK(clk), .RN(n529), .Q(
        \CACHE[1][107] ), .QN(n803) );
  DFFRX1 \CACHE_reg[1][106]  ( .D(n2042), .CK(clk), .RN(n531), .Q(
        \CACHE[1][106] ), .QN(n802) );
  DFFRX1 \CACHE_reg[1][105]  ( .D(n2041), .CK(clk), .RN(n534), .Q(
        \CACHE[1][105] ), .QN(n801) );
  DFFRX1 \CACHE_reg[1][104]  ( .D(n2040), .CK(clk), .RN(n537), .Q(
        \CACHE[1][104] ), .QN(n800) );
  DFFRX1 \CACHE_reg[1][103]  ( .D(n2039), .CK(clk), .RN(n539), .Q(
        \CACHE[1][103] ), .QN(n799) );
  DFFRX1 \CACHE_reg[1][102]  ( .D(n2038), .CK(clk), .RN(n3022), .Q(
        \CACHE[1][102] ), .QN(n798) );
  DFFRX1 \CACHE_reg[1][101]  ( .D(n2037), .CK(clk), .RN(n3025), .Q(
        \CACHE[1][101] ), .QN(n797) );
  DFFRX1 \CACHE_reg[1][100]  ( .D(n2036), .CK(clk), .RN(n3034), .Q(
        \CACHE[1][100] ), .QN(n796) );
  DFFRX1 \CACHE_reg[1][99]  ( .D(n2035), .CK(clk), .RN(n3027), .Q(
        \CACHE[1][99] ), .QN(n795) );
  DFFRX1 \CACHE_reg[1][98]  ( .D(n2034), .CK(clk), .RN(n3030), .Q(
        \CACHE[1][98] ), .QN(n794) );
  DFFRX1 \CACHE_reg[1][97]  ( .D(n2033), .CK(clk), .RN(n3035), .Q(
        \CACHE[1][97] ), .QN(n793) );
  DFFRX1 \CACHE_reg[1][96]  ( .D(n2032), .CK(clk), .RN(n3033), .Q(
        \CACHE[1][96] ), .QN(n792) );
  DFFRX1 \CACHE_reg[1][95]  ( .D(n2031), .CK(clk), .RN(n477), .Q(
        \CACHE[1][95] ), .QN(n791) );
  DFFRX1 \CACHE_reg[1][94]  ( .D(n2030), .CK(clk), .RN(n480), .Q(
        \CACHE[1][94] ), .QN(n790) );
  DFFRX1 \CACHE_reg[1][93]  ( .D(n2029), .CK(clk), .RN(n483), .Q(
        \CACHE[1][93] ), .QN(n789) );
  DFFRX1 \CACHE_reg[1][92]  ( .D(n2028), .CK(clk), .RN(n485), .Q(
        \CACHE[1][92] ), .QN(n788) );
  DFFRX1 \CACHE_reg[1][91]  ( .D(n2027), .CK(clk), .RN(n488), .Q(
        \CACHE[1][91] ), .QN(n787) );
  DFFRX1 \CACHE_reg[1][90]  ( .D(n2026), .CK(clk), .RN(n491), .Q(
        \CACHE[1][90] ), .QN(n786) );
  DFFRX1 \CACHE_reg[1][89]  ( .D(n2025), .CK(clk), .RN(n493), .Q(
        \CACHE[1][89] ), .QN(n785) );
  DFFRX1 \CACHE_reg[1][88]  ( .D(n2024), .CK(clk), .RN(n496), .Q(
        \CACHE[1][88] ), .QN(n784) );
  DFFRX1 \CACHE_reg[1][87]  ( .D(n2023), .CK(clk), .RN(n499), .Q(
        \CACHE[1][87] ), .QN(n783) );
  DFFRX1 \CACHE_reg[1][86]  ( .D(n2022), .CK(clk), .RN(n501), .Q(
        \CACHE[1][86] ), .QN(n782) );
  DFFRX1 \CACHE_reg[1][85]  ( .D(n2021), .CK(clk), .RN(n504), .Q(
        \CACHE[1][85] ), .QN(n781) );
  DFFRX1 \CACHE_reg[1][84]  ( .D(n2020), .CK(clk), .RN(n507), .Q(
        \CACHE[1][84] ), .QN(n780) );
  DFFRX1 \CACHE_reg[1][83]  ( .D(n2019), .CK(clk), .RN(n509), .Q(
        \CACHE[1][83] ), .QN(n779) );
  DFFRX1 \CACHE_reg[1][82]  ( .D(n2018), .CK(clk), .RN(n3035), .Q(
        \CACHE[1][82] ), .QN(n778) );
  DFFRX1 \CACHE_reg[1][81]  ( .D(n2017), .CK(clk), .RN(n512), .Q(
        \CACHE[1][81] ), .QN(n777) );
  DFFRX1 \CACHE_reg[1][80]  ( .D(n2016), .CK(clk), .RN(n515), .Q(
        \CACHE[1][80] ), .QN(n776) );
  DFFRX1 \CACHE_reg[1][79]  ( .D(n2015), .CK(clk), .RN(n517), .Q(
        \CACHE[1][79] ), .QN(n775) );
  DFFRX1 \CACHE_reg[1][78]  ( .D(n2014), .CK(clk), .RN(n520), .Q(
        \CACHE[1][78] ), .QN(n774) );
  DFFRX1 \CACHE_reg[1][77]  ( .D(n2013), .CK(clk), .RN(n523), .Q(
        \CACHE[1][77] ), .QN(n773) );
  DFFRX1 \CACHE_reg[1][76]  ( .D(n2012), .CK(clk), .RN(n525), .Q(
        \CACHE[1][76] ), .QN(n772) );
  DFFRX1 \CACHE_reg[1][75]  ( .D(n2011), .CK(clk), .RN(n528), .Q(
        \CACHE[1][75] ), .QN(n771) );
  DFFRX1 \CACHE_reg[1][74]  ( .D(n2010), .CK(clk), .RN(n531), .Q(
        \CACHE[1][74] ), .QN(n770) );
  DFFRX1 \CACHE_reg[1][73]  ( .D(n2009), .CK(clk), .RN(n533), .Q(
        \CACHE[1][73] ), .QN(n769) );
  DFFRX1 \CACHE_reg[1][72]  ( .D(n2008), .CK(clk), .RN(n536), .Q(
        \CACHE[1][72] ), .QN(n768) );
  DFFRX1 \CACHE_reg[1][71]  ( .D(n2007), .CK(clk), .RN(n539), .Q(
        \CACHE[1][71] ), .QN(n767) );
  DFFRX1 \CACHE_reg[1][70]  ( .D(n2006), .CK(clk), .RN(n3020), .Q(
        \CACHE[1][70] ), .QN(n766) );
  DFFRX1 \CACHE_reg[1][69]  ( .D(n2005), .CK(clk), .RN(n3024), .Q(
        \CACHE[1][69] ), .QN(n765) );
  DFFRX1 \CACHE_reg[1][68]  ( .D(n2004), .CK(clk), .RN(n3036), .Q(
        \CACHE[1][68] ), .QN(n764) );
  DFFRX1 \CACHE_reg[1][67]  ( .D(n2003), .CK(clk), .RN(n3027), .Q(
        \CACHE[1][67] ), .QN(n763) );
  DFFRX1 \CACHE_reg[1][66]  ( .D(n2002), .CK(clk), .RN(n3029), .Q(
        \CACHE[1][66] ), .QN(n762) );
  DFFRX1 \CACHE_reg[1][65]  ( .D(n2001), .CK(clk), .RN(n3037), .Q(
        \CACHE[1][65] ), .QN(n761) );
  DFFRX1 \CACHE_reg[1][64]  ( .D(n2000), .CK(clk), .RN(n3032), .Q(
        \CACHE[1][64] ), .QN(n760) );
  DFFRX1 \CACHE_reg[1][63]  ( .D(n1999), .CK(clk), .RN(n477), .Q(
        \CACHE[1][63] ), .QN(n759) );
  DFFRX1 \CACHE_reg[1][62]  ( .D(n1998), .CK(clk), .RN(n479), .Q(
        \CACHE[1][62] ), .QN(n758) );
  DFFRX1 \CACHE_reg[1][61]  ( .D(n1997), .CK(clk), .RN(n482), .Q(
        \CACHE[1][61] ), .QN(n757) );
  DFFRX1 \CACHE_reg[1][60]  ( .D(n1996), .CK(clk), .RN(n485), .Q(
        \CACHE[1][60] ), .QN(n756) );
  DFFRX1 \CACHE_reg[1][59]  ( .D(n1995), .CK(clk), .RN(n487), .Q(
        \CACHE[1][59] ), .QN(n755) );
  DFFRX1 \CACHE_reg[1][58]  ( .D(n1994), .CK(clk), .RN(n490), .Q(
        \CACHE[1][58] ), .QN(n754) );
  DFFRX1 \CACHE_reg[1][57]  ( .D(n1993), .CK(clk), .RN(n493), .Q(
        \CACHE[1][57] ), .QN(n753) );
  DFFRX1 \CACHE_reg[1][56]  ( .D(n1992), .CK(clk), .RN(n495), .Q(
        \CACHE[1][56] ), .QN(n752) );
  DFFRX1 \CACHE_reg[1][55]  ( .D(n1991), .CK(clk), .RN(n498), .Q(
        \CACHE[1][55] ), .QN(n751) );
  DFFRX1 \CACHE_reg[1][54]  ( .D(n1990), .CK(clk), .RN(n501), .Q(
        \CACHE[1][54] ), .QN(n750) );
  DFFRX1 \CACHE_reg[1][53]  ( .D(n1989), .CK(clk), .RN(n503), .Q(
        \CACHE[1][53] ), .QN(n749) );
  DFFRX1 \CACHE_reg[1][52]  ( .D(n1988), .CK(clk), .RN(n506), .Q(
        \CACHE[1][52] ), .QN(n748) );
  DFFRX1 \CACHE_reg[1][51]  ( .D(n1987), .CK(clk), .RN(n509), .Q(
        \CACHE[1][51] ), .QN(n747) );
  DFFRX1 \CACHE_reg[1][50]  ( .D(n1986), .CK(clk), .RN(n3037), .Q(
        \CACHE[1][50] ), .QN(n746) );
  DFFRX1 \CACHE_reg[1][49]  ( .D(n1985), .CK(clk), .RN(n511), .Q(
        \CACHE[1][49] ), .QN(n745) );
  DFFRX1 \CACHE_reg[1][48]  ( .D(n1984), .CK(clk), .RN(n514), .Q(
        \CACHE[1][48] ), .QN(n744) );
  DFFRX1 \CACHE_reg[1][47]  ( .D(n1983), .CK(clk), .RN(n517), .Q(
        \CACHE[1][47] ), .QN(n743) );
  DFFRX1 \CACHE_reg[1][46]  ( .D(n1982), .CK(clk), .RN(n519), .Q(
        \CACHE[1][46] ), .QN(n742) );
  DFFRX1 \CACHE_reg[1][45]  ( .D(n1981), .CK(clk), .RN(n522), .Q(
        \CACHE[1][45] ), .QN(n741) );
  DFFRX1 \CACHE_reg[1][44]  ( .D(n1980), .CK(clk), .RN(n525), .Q(
        \CACHE[1][44] ), .QN(n740) );
  DFFRX1 \CACHE_reg[1][43]  ( .D(n1979), .CK(clk), .RN(n527), .Q(
        \CACHE[1][43] ), .QN(n739) );
  DFFRX1 \CACHE_reg[1][42]  ( .D(n1978), .CK(clk), .RN(n530), .Q(
        \CACHE[1][42] ), .QN(n738) );
  DFFRX1 \CACHE_reg[1][41]  ( .D(n1977), .CK(clk), .RN(n533), .Q(
        \CACHE[1][41] ), .QN(n737) );
  DFFRX1 \CACHE_reg[1][40]  ( .D(n1976), .CK(clk), .RN(n535), .Q(
        \CACHE[1][40] ), .QN(n736) );
  DFFRX1 \CACHE_reg[1][39]  ( .D(n1975), .CK(clk), .RN(n538), .Q(
        \CACHE[1][39] ), .QN(n735) );
  DFFRX1 \CACHE_reg[1][38]  ( .D(n1974), .CK(clk), .RN(n3020), .Q(
        \CACHE[1][38] ), .QN(n734) );
  DFFRX1 \CACHE_reg[1][37]  ( .D(n1973), .CK(clk), .RN(n3023), .Q(
        \CACHE[1][37] ), .QN(n733) );
  DFFRX1 \CACHE_reg[1][36]  ( .D(n1972), .CK(clk), .RN(n3038), .Q(
        \CACHE[1][36] ), .QN(n732) );
  DFFRX1 \CACHE_reg[1][35]  ( .D(n1971), .CK(clk), .RN(n3026), .Q(
        \CACHE[1][35] ), .QN(n731) );
  DFFRX1 \CACHE_reg[1][34]  ( .D(n1970), .CK(clk), .RN(n3029), .Q(
        \CACHE[1][34] ), .QN(n730) );
  DFFRX1 \CACHE_reg[1][33]  ( .D(n1969), .CK(clk), .RN(n3039), .Q(
        \CACHE[1][33] ), .QN(n729) );
  DFFRX1 \CACHE_reg[1][32]  ( .D(n1968), .CK(clk), .RN(n3031), .Q(
        \CACHE[1][32] ), .QN(n728) );
  DFFRX1 \CACHE_reg[1][31]  ( .D(n1967), .CK(clk), .RN(n476), .Q(
        \CACHE[1][31] ), .QN(n727) );
  DFFRX1 \CACHE_reg[1][30]  ( .D(n1966), .CK(clk), .RN(n479), .Q(
        \CACHE[1][30] ), .QN(n726) );
  DFFRX1 \CACHE_reg[1][29]  ( .D(n1965), .CK(clk), .RN(n481), .Q(
        \CACHE[1][29] ), .QN(n725) );
  DFFRX1 \CACHE_reg[1][28]  ( .D(n1964), .CK(clk), .RN(n484), .Q(
        \CACHE[1][28] ), .QN(n724) );
  DFFRX1 \CACHE_reg[1][27]  ( .D(n1963), .CK(clk), .RN(n487), .Q(
        \CACHE[1][27] ), .QN(n723) );
  DFFRX1 \CACHE_reg[1][26]  ( .D(n1962), .CK(clk), .RN(n489), .Q(
        \CACHE[1][26] ), .QN(n722) );
  DFFRX1 \CACHE_reg[1][25]  ( .D(n1961), .CK(clk), .RN(n492), .Q(
        \CACHE[1][25] ), .QN(n721) );
  DFFRX1 \CACHE_reg[1][24]  ( .D(n1960), .CK(clk), .RN(n495), .Q(
        \CACHE[1][24] ), .QN(n720) );
  DFFRX1 \CACHE_reg[1][23]  ( .D(n1959), .CK(clk), .RN(n497), .Q(
        \CACHE[1][23] ), .QN(n719) );
  DFFRX1 \CACHE_reg[1][22]  ( .D(n1958), .CK(clk), .RN(n500), .Q(
        \CACHE[1][22] ), .QN(n718) );
  DFFRX1 \CACHE_reg[1][21]  ( .D(n1957), .CK(clk), .RN(n503), .Q(
        \CACHE[1][21] ), .QN(n717) );
  DFFRX1 \CACHE_reg[1][20]  ( .D(n1956), .CK(clk), .RN(n505), .Q(
        \CACHE[1][20] ), .QN(n716) );
  DFFRX1 \CACHE_reg[1][19]  ( .D(n1955), .CK(clk), .RN(n508), .Q(
        \CACHE[1][19] ), .QN(n715) );
  DFFRX1 \CACHE_reg[1][18]  ( .D(n1954), .CK(clk), .RN(n3059), .Q(
        \CACHE[1][18] ), .QN(n714) );
  DFFRX1 \CACHE_reg[1][17]  ( .D(n1953), .CK(clk), .RN(n511), .Q(
        \CACHE[1][17] ), .QN(n713) );
  DFFRX1 \CACHE_reg[1][16]  ( .D(n1952), .CK(clk), .RN(n513), .Q(
        \CACHE[1][16] ), .QN(n712) );
  DFFRX1 \CACHE_reg[1][15]  ( .D(n1951), .CK(clk), .RN(n516), .Q(
        \CACHE[1][15] ), .QN(n711) );
  DFFRX1 \CACHE_reg[1][14]  ( .D(n1950), .CK(clk), .RN(n519), .Q(
        \CACHE[1][14] ), .QN(n710) );
  DFFRX1 \CACHE_reg[1][13]  ( .D(n1949), .CK(clk), .RN(n521), .Q(
        \CACHE[1][13] ), .QN(n709) );
  DFFRX1 \CACHE_reg[1][12]  ( .D(n1948), .CK(clk), .RN(n524), .Q(
        \CACHE[1][12] ), .QN(n708) );
  DFFRX1 \CACHE_reg[1][11]  ( .D(n1947), .CK(clk), .RN(n527), .Q(
        \CACHE[1][11] ), .QN(n707) );
  DFFRX1 \CACHE_reg[1][10]  ( .D(n1946), .CK(clk), .RN(n529), .Q(
        \CACHE[1][10] ), .QN(n706) );
  DFFRX1 \CACHE_reg[1][9]  ( .D(n1945), .CK(clk), .RN(n532), .Q(\CACHE[1][9] ), 
        .QN(n705) );
  DFFRX1 \CACHE_reg[1][8]  ( .D(n1944), .CK(clk), .RN(n535), .Q(\CACHE[1][8] ), 
        .QN(n704) );
  DFFRX1 \CACHE_reg[1][7]  ( .D(n1943), .CK(clk), .RN(n537), .Q(\CACHE[1][7] ), 
        .QN(n703) );
  DFFRX1 \CACHE_reg[1][6]  ( .D(n1942), .CK(clk), .RN(n540), .Q(\CACHE[1][6] ), 
        .QN(n702) );
  DFFRX1 \CACHE_reg[1][5]  ( .D(n1941), .CK(clk), .RN(n3023), .Q(\CACHE[1][5] ), .QN(n701) );
  DFFRX1 \CACHE_reg[1][4]  ( .D(n1940), .CK(clk), .RN(n3058), .Q(\CACHE[1][4] ), .QN(n700) );
  DFFRX1 \CACHE_reg[1][3]  ( .D(n1939), .CK(clk), .RN(n3025), .Q(\CACHE[1][3] ), .QN(n699) );
  DFFRX1 \CACHE_reg[1][2]  ( .D(n1938), .CK(clk), .RN(n3028), .Q(\CACHE[1][2] ), .QN(n698) );
  DFFRX1 \CACHE_reg[1][1]  ( .D(n1937), .CK(clk), .RN(n3039), .Q(\CACHE[1][1] ), .QN(n697) );
  DFFRX1 \CACHE_reg[1][0]  ( .D(n1936), .CK(clk), .RN(n3031), .Q(\CACHE[1][0] ), .QN(n696) );
  DFFRX1 \CACHE_reg[4][154]  ( .D(n2555), .CK(clk), .RN(n3057), .Q(
        \CACHE[4][154] ), .QN(n1315) );
  DFFRX1 \CACHE_reg[4][153]  ( .D(n2554), .CK(clk), .RN(n3056), .Q(
        \CACHE[4][153] ), .QN(n1314) );
  DFFRX1 \CACHE_reg[4][152]  ( .D(n2553), .CK(clk), .RN(n3056), .Q(
        \CACHE[4][152] ), .QN(n1313) );
  DFFRX1 \CACHE_reg[4][151]  ( .D(n2552), .CK(clk), .RN(n3040), .Q(
        \CACHE[4][151] ), .QN(n1312) );
  DFFRX1 \CACHE_reg[4][150]  ( .D(n2551), .CK(clk), .RN(n3040), .Q(
        \CACHE[4][150] ), .QN(n1311) );
  DFFRX1 \CACHE_reg[4][149]  ( .D(n2550), .CK(clk), .RN(n3041), .Q(
        \CACHE[4][149] ), .QN(n1310) );
  DFFRX1 \CACHE_reg[4][148]  ( .D(n2549), .CK(clk), .RN(n3042), .Q(
        \CACHE[4][148] ), .QN(n1309) );
  DFFRX1 \CACHE_reg[4][147]  ( .D(n2548), .CK(clk), .RN(n3042), .Q(
        \CACHE[4][147] ), .QN(n1308) );
  DFFRX1 \CACHE_reg[4][146]  ( .D(n2547), .CK(clk), .RN(n3043), .Q(
        \CACHE[4][146] ), .QN(n1307) );
  DFFRX1 \CACHE_reg[4][145]  ( .D(n2546), .CK(clk), .RN(n3044), .Q(
        \CACHE[4][145] ), .QN(n1306) );
  DFFRX1 \CACHE_reg[4][144]  ( .D(n2545), .CK(clk), .RN(n3044), .Q(
        \CACHE[4][144] ), .QN(n1305) );
  DFFRX1 \CACHE_reg[4][143]  ( .D(n2544), .CK(clk), .RN(n3045), .Q(
        \CACHE[4][143] ), .QN(n1304) );
  DFFRX1 \CACHE_reg[4][142]  ( .D(n2543), .CK(clk), .RN(n3046), .Q(
        \CACHE[4][142] ), .QN(n1303) );
  DFFRX1 \CACHE_reg[4][141]  ( .D(n2542), .CK(clk), .RN(n3046), .Q(
        \CACHE[4][141] ), .QN(n1302) );
  DFFRX1 \CACHE_reg[4][140]  ( .D(n2541), .CK(clk), .RN(n3047), .Q(
        \CACHE[4][140] ), .QN(n1301) );
  DFFRX1 \CACHE_reg[4][139]  ( .D(n2540), .CK(clk), .RN(n3048), .Q(
        \CACHE[4][139] ), .QN(n1300) );
  DFFRX1 \CACHE_reg[4][138]  ( .D(n2539), .CK(clk), .RN(n3048), .Q(
        \CACHE[4][138] ), .QN(n1299) );
  DFFRX1 \CACHE_reg[4][137]  ( .D(n2538), .CK(clk), .RN(n3049), .Q(
        \CACHE[4][137] ), .QN(n1298) );
  DFFRX1 \CACHE_reg[4][136]  ( .D(n2537), .CK(clk), .RN(n3050), .Q(
        \CACHE[4][136] ), .QN(n1297) );
  DFFRX1 \CACHE_reg[4][135]  ( .D(n2536), .CK(clk), .RN(n3050), .Q(
        \CACHE[4][135] ), .QN(n1296) );
  DFFRX1 \CACHE_reg[4][134]  ( .D(n2535), .CK(clk), .RN(n3051), .Q(
        \CACHE[4][134] ), .QN(n1295) );
  DFFRX1 \CACHE_reg[4][133]  ( .D(n2534), .CK(clk), .RN(n3052), .Q(
        \CACHE[4][133] ), .QN(n1294) );
  DFFRX1 \CACHE_reg[4][132]  ( .D(n2533), .CK(clk), .RN(n3052), .Q(
        \CACHE[4][132] ), .QN(n1293) );
  DFFRX1 \CACHE_reg[4][131]  ( .D(n2532), .CK(clk), .RN(n3053), .Q(
        \CACHE[4][131] ), .QN(n1292) );
  DFFRX1 \CACHE_reg[4][130]  ( .D(n2531), .CK(clk), .RN(n3054), .Q(
        \CACHE[4][130] ), .QN(n1291) );
  DFFRX1 \CACHE_reg[4][129]  ( .D(n2530), .CK(clk), .RN(n3054), .Q(
        \CACHE[4][129] ), .QN(n1290) );
  DFFRX1 \CACHE_reg[4][128]  ( .D(n2529), .CK(clk), .RN(n3055), .Q(
        \CACHE[4][128] ), .QN(n1289) );
  DFFRX1 \CACHE_reg[4][127]  ( .D(n2528), .CK(clk), .RN(n478), .Q(
        \CACHE[4][127] ), .QN(n1288) );
  DFFRX1 \CACHE_reg[4][126]  ( .D(n2527), .CK(clk), .RN(n480), .Q(
        \CACHE[4][126] ), .QN(n1287) );
  DFFRX1 \CACHE_reg[4][125]  ( .D(n2526), .CK(clk), .RN(n483), .Q(
        \CACHE[4][125] ), .QN(n1286) );
  DFFRX1 \CACHE_reg[4][124]  ( .D(n2525), .CK(clk), .RN(n486), .Q(
        \CACHE[4][124] ), .QN(n1285) );
  DFFRX1 \CACHE_reg[4][123]  ( .D(n2524), .CK(clk), .RN(n488), .Q(
        \CACHE[4][123] ), .QN(n1284) );
  DFFRX1 \CACHE_reg[4][122]  ( .D(n2523), .CK(clk), .RN(n491), .Q(
        \CACHE[4][122] ), .QN(n1283) );
  DFFRX1 \CACHE_reg[4][121]  ( .D(n2522), .CK(clk), .RN(n494), .Q(
        \CACHE[4][121] ), .QN(n1282) );
  DFFRX1 \CACHE_reg[4][120]  ( .D(n2521), .CK(clk), .RN(n496), .Q(
        \CACHE[4][120] ), .QN(n1281) );
  DFFRX1 \CACHE_reg[4][119]  ( .D(n2520), .CK(clk), .RN(n499), .Q(
        \CACHE[4][119] ), .QN(n1280) );
  DFFRX1 \CACHE_reg[4][118]  ( .D(n2519), .CK(clk), .RN(n502), .Q(
        \CACHE[4][118] ), .QN(n1279) );
  DFFRX1 \CACHE_reg[4][117]  ( .D(n2518), .CK(clk), .RN(n504), .Q(
        \CACHE[4][117] ), .QN(n1278) );
  DFFRX1 \CACHE_reg[4][116]  ( .D(n2517), .CK(clk), .RN(n507), .Q(
        \CACHE[4][116] ), .QN(n1277) );
  DFFRX1 \CACHE_reg[4][115]  ( .D(n2516), .CK(clk), .RN(n510), .Q(
        \CACHE[4][115] ), .QN(n1276) );
  DFFRX1 \CACHE_reg[4][114]  ( .D(n2515), .CK(clk), .RN(n3033), .Q(
        \CACHE[4][114] ), .QN(n1275) );
  DFFRX1 \CACHE_reg[4][113]  ( .D(n2514), .CK(clk), .RN(n512), .Q(
        \CACHE[4][113] ), .QN(n1274) );
  DFFRX1 \CACHE_reg[4][112]  ( .D(n2513), .CK(clk), .RN(n515), .Q(
        \CACHE[4][112] ), .QN(n1273) );
  DFFRX1 \CACHE_reg[4][111]  ( .D(n2512), .CK(clk), .RN(n518), .Q(
        \CACHE[4][111] ), .QN(n1272) );
  DFFRX1 \CACHE_reg[4][110]  ( .D(n2511), .CK(clk), .RN(n520), .Q(
        \CACHE[4][110] ), .QN(n1271) );
  DFFRX1 \CACHE_reg[4][109]  ( .D(n2510), .CK(clk), .RN(n523), .Q(
        \CACHE[4][109] ), .QN(n1270) );
  DFFRX1 \CACHE_reg[4][108]  ( .D(n2509), .CK(clk), .RN(n526), .Q(
        \CACHE[4][108] ), .QN(n1269) );
  DFFRX1 \CACHE_reg[4][107]  ( .D(n2508), .CK(clk), .RN(n528), .Q(
        \CACHE[4][107] ), .QN(n1268) );
  DFFRX1 \CACHE_reg[4][106]  ( .D(n2507), .CK(clk), .RN(n531), .Q(
        \CACHE[4][106] ), .QN(n1267) );
  DFFRX1 \CACHE_reg[4][105]  ( .D(n2506), .CK(clk), .RN(n534), .Q(
        \CACHE[4][105] ), .QN(n1266) );
  DFFRX1 \CACHE_reg[4][104]  ( .D(n2505), .CK(clk), .RN(n536), .Q(
        \CACHE[4][104] ), .QN(n1265) );
  DFFRX1 \CACHE_reg[4][103]  ( .D(n2504), .CK(clk), .RN(n539), .Q(
        \CACHE[4][103] ), .QN(n1264) );
  DFFRX1 \CACHE_reg[4][102]  ( .D(n2503), .CK(clk), .RN(n3022), .Q(
        \CACHE[4][102] ), .QN(n1263) );
  DFFRX1 \CACHE_reg[4][101]  ( .D(n2502), .CK(clk), .RN(n3024), .Q(
        \CACHE[4][101] ), .QN(n1262) );
  DFFRX1 \CACHE_reg[4][100]  ( .D(n2501), .CK(clk), .RN(n3034), .Q(
        \CACHE[4][100] ), .QN(n1261) );
  DFFRX1 \CACHE_reg[4][99]  ( .D(n2500), .CK(clk), .RN(n3027), .Q(
        \CACHE[4][99] ), .QN(n1260) );
  DFFRX1 \CACHE_reg[4][98]  ( .D(n2499), .CK(clk), .RN(n3030), .Q(
        \CACHE[4][98] ), .QN(n1259) );
  DFFRX1 \CACHE_reg[4][97]  ( .D(n2498), .CK(clk), .RN(n3034), .Q(
        \CACHE[4][97] ), .QN(n1258) );
  DFFRX1 \CACHE_reg[4][96]  ( .D(n2497), .CK(clk), .RN(n3032), .Q(
        \CACHE[4][96] ), .QN(n1257) );
  DFFRX1 \CACHE_reg[4][95]  ( .D(n2496), .CK(clk), .RN(n477), .Q(
        \CACHE[4][95] ), .QN(n1256) );
  DFFRX1 \CACHE_reg[4][94]  ( .D(n2495), .CK(clk), .RN(n480), .Q(
        \CACHE[4][94] ), .QN(n1255) );
  DFFRX1 \CACHE_reg[4][93]  ( .D(n2494), .CK(clk), .RN(n482), .Q(
        \CACHE[4][93] ), .QN(n1254) );
  DFFRX1 \CACHE_reg[4][92]  ( .D(n2493), .CK(clk), .RN(n485), .Q(
        \CACHE[4][92] ), .QN(n1253) );
  DFFRX1 \CACHE_reg[4][91]  ( .D(n2492), .CK(clk), .RN(n488), .Q(
        \CACHE[4][91] ), .QN(n1252) );
  DFFRX1 \CACHE_reg[4][90]  ( .D(n2491), .CK(clk), .RN(n490), .Q(
        \CACHE[4][90] ), .QN(n1251) );
  DFFRX1 \CACHE_reg[4][89]  ( .D(n2490), .CK(clk), .RN(n493), .Q(
        \CACHE[4][89] ), .QN(n1250) );
  DFFRX1 \CACHE_reg[4][88]  ( .D(n2489), .CK(clk), .RN(n496), .Q(
        \CACHE[4][88] ), .QN(n1249) );
  DFFRX1 \CACHE_reg[4][87]  ( .D(n2488), .CK(clk), .RN(n498), .Q(
        \CACHE[4][87] ), .QN(n1248) );
  DFFRX1 \CACHE_reg[4][86]  ( .D(n2487), .CK(clk), .RN(n501), .Q(
        \CACHE[4][86] ), .QN(n1247) );
  DFFRX1 \CACHE_reg[4][85]  ( .D(n2486), .CK(clk), .RN(n504), .Q(
        \CACHE[4][85] ), .QN(n1246) );
  DFFRX1 \CACHE_reg[4][84]  ( .D(n2485), .CK(clk), .RN(n506), .Q(
        \CACHE[4][84] ), .QN(n1245) );
  DFFRX1 \CACHE_reg[4][83]  ( .D(n2484), .CK(clk), .RN(n509), .Q(
        \CACHE[4][83] ), .QN(n1244) );
  DFFRX1 \CACHE_reg[4][82]  ( .D(n2483), .CK(clk), .RN(n3035), .Q(
        \CACHE[4][82] ), .QN(n1243) );
  DFFRX1 \CACHE_reg[4][81]  ( .D(n2482), .CK(clk), .RN(n512), .Q(
        \CACHE[4][81] ), .QN(n1242) );
  DFFRX1 \CACHE_reg[4][80]  ( .D(n2481), .CK(clk), .RN(n514), .Q(
        \CACHE[4][80] ), .QN(n1241) );
  DFFRX1 \CACHE_reg[4][79]  ( .D(n2480), .CK(clk), .RN(n517), .Q(
        \CACHE[4][79] ), .QN(n1240) );
  DFFRX1 \CACHE_reg[4][78]  ( .D(n2479), .CK(clk), .RN(n520), .Q(
        \CACHE[4][78] ), .QN(n1239) );
  DFFRX1 \CACHE_reg[4][77]  ( .D(n2478), .CK(clk), .RN(n522), .Q(
        \CACHE[4][77] ), .QN(n1238) );
  DFFRX1 \CACHE_reg[4][76]  ( .D(n2477), .CK(clk), .RN(n525), .Q(
        \CACHE[4][76] ), .QN(n1237) );
  DFFRX1 \CACHE_reg[4][75]  ( .D(n2476), .CK(clk), .RN(n528), .Q(
        \CACHE[4][75] ), .QN(n1236) );
  DFFRX1 \CACHE_reg[4][74]  ( .D(n2475), .CK(clk), .RN(n530), .Q(
        \CACHE[4][74] ), .QN(n1235) );
  DFFRX1 \CACHE_reg[4][73]  ( .D(n2474), .CK(clk), .RN(n533), .Q(
        \CACHE[4][73] ), .QN(n1234) );
  DFFRX1 \CACHE_reg[4][72]  ( .D(n2473), .CK(clk), .RN(n536), .Q(
        \CACHE[4][72] ), .QN(n1233) );
  DFFRX1 \CACHE_reg[4][71]  ( .D(n2472), .CK(clk), .RN(n538), .Q(
        \CACHE[4][71] ), .QN(n1232) );
  DFFRX1 \CACHE_reg[4][70]  ( .D(n2471), .CK(clk), .RN(n3020), .Q(
        \CACHE[4][70] ), .QN(n1231) );
  DFFRX1 \CACHE_reg[4][69]  ( .D(n2470), .CK(clk), .RN(n3024), .Q(
        \CACHE[4][69] ), .QN(n1230) );
  DFFRX1 \CACHE_reg[4][68]  ( .D(n2469), .CK(clk), .RN(n3036), .Q(
        \CACHE[4][68] ), .QN(n1229) );
  DFFRX1 \CACHE_reg[4][67]  ( .D(n2468), .CK(clk), .RN(n3026), .Q(
        \CACHE[4][67] ), .QN(n1228) );
  DFFRX1 \CACHE_reg[4][66]  ( .D(n2467), .CK(clk), .RN(n3029), .Q(
        \CACHE[4][66] ), .QN(n1227) );
  DFFRX1 \CACHE_reg[4][65]  ( .D(n2466), .CK(clk), .RN(n3036), .Q(
        \CACHE[4][65] ), .QN(n1226) );
  DFFRX1 \CACHE_reg[4][64]  ( .D(n2465), .CK(clk), .RN(n3032), .Q(
        \CACHE[4][64] ), .QN(n1225) );
  DFFRX1 \CACHE_reg[4][63]  ( .D(n2464), .CK(clk), .RN(n476), .Q(
        \CACHE[4][63] ), .QN(n1224) );
  DFFRX1 \CACHE_reg[4][62]  ( .D(n2463), .CK(clk), .RN(n479), .Q(
        \CACHE[4][62] ), .QN(n1223) );
  DFFRX1 \CACHE_reg[4][61]  ( .D(n2462), .CK(clk), .RN(n482), .Q(
        \CACHE[4][61] ), .QN(n1222) );
  DFFRX1 \CACHE_reg[4][60]  ( .D(n2461), .CK(clk), .RN(n484), .Q(
        \CACHE[4][60] ), .QN(n1221) );
  DFFRX1 \CACHE_reg[4][59]  ( .D(n2460), .CK(clk), .RN(n487), .Q(
        \CACHE[4][59] ), .QN(n1220) );
  DFFRX1 \CACHE_reg[4][58]  ( .D(n2459), .CK(clk), .RN(n490), .Q(
        \CACHE[4][58] ), .QN(n1219) );
  DFFRX1 \CACHE_reg[4][57]  ( .D(n2458), .CK(clk), .RN(n492), .Q(
        \CACHE[4][57] ), .QN(n1218) );
  DFFRX1 \CACHE_reg[4][56]  ( .D(n2457), .CK(clk), .RN(n495), .Q(
        \CACHE[4][56] ), .QN(n1217) );
  DFFRX1 \CACHE_reg[4][55]  ( .D(n2456), .CK(clk), .RN(n498), .Q(
        \CACHE[4][55] ), .QN(n1216) );
  DFFRX1 \CACHE_reg[4][54]  ( .D(n2455), .CK(clk), .RN(n500), .Q(
        \CACHE[4][54] ), .QN(n1215) );
  DFFRX1 \CACHE_reg[4][53]  ( .D(n2454), .CK(clk), .RN(n503), .Q(
        \CACHE[4][53] ), .QN(n1214) );
  DFFRX1 \CACHE_reg[4][52]  ( .D(n2453), .CK(clk), .RN(n506), .Q(
        \CACHE[4][52] ), .QN(n1213) );
  DFFRX1 \CACHE_reg[4][51]  ( .D(n2452), .CK(clk), .RN(n508), .Q(
        \CACHE[4][51] ), .QN(n1212) );
  DFFRX1 \CACHE_reg[4][50]  ( .D(n2451), .CK(clk), .RN(n3037), .Q(
        \CACHE[4][50] ), .QN(n1211) );
  DFFRX1 \CACHE_reg[4][49]  ( .D(n2450), .CK(clk), .RN(n511), .Q(
        \CACHE[4][49] ), .QN(n1210) );
  DFFRX1 \CACHE_reg[4][48]  ( .D(n2449), .CK(clk), .RN(n514), .Q(
        \CACHE[4][48] ), .QN(n1209) );
  DFFRX1 \CACHE_reg[4][47]  ( .D(n2448), .CK(clk), .RN(n516), .Q(
        \CACHE[4][47] ), .QN(n1208) );
  DFFRX1 \CACHE_reg[4][46]  ( .D(n2447), .CK(clk), .RN(n519), .Q(
        \CACHE[4][46] ), .QN(n1207) );
  DFFRX1 \CACHE_reg[4][45]  ( .D(n2446), .CK(clk), .RN(n522), .Q(
        \CACHE[4][45] ), .QN(n1206) );
  DFFRX1 \CACHE_reg[4][44]  ( .D(n2445), .CK(clk), .RN(n524), .Q(
        \CACHE[4][44] ), .QN(n1205) );
  DFFRX1 \CACHE_reg[4][43]  ( .D(n2444), .CK(clk), .RN(n527), .Q(
        \CACHE[4][43] ), .QN(n1204) );
  DFFRX1 \CACHE_reg[4][42]  ( .D(n2443), .CK(clk), .RN(n530), .Q(
        \CACHE[4][42] ), .QN(n1203) );
  DFFRX1 \CACHE_reg[4][41]  ( .D(n2442), .CK(clk), .RN(n532), .Q(
        \CACHE[4][41] ), .QN(n1202) );
  DFFRX1 \CACHE_reg[4][40]  ( .D(n2441), .CK(clk), .RN(n535), .Q(
        \CACHE[4][40] ), .QN(n1201) );
  DFFRX1 \CACHE_reg[4][39]  ( .D(n2440), .CK(clk), .RN(n538), .Q(
        \CACHE[4][39] ), .QN(n1200) );
  DFFRX1 \CACHE_reg[4][38]  ( .D(n2439), .CK(clk), .RN(n540), .Q(
        \CACHE[4][38] ), .QN(n1199) );
  DFFRX1 \CACHE_reg[4][37]  ( .D(n2438), .CK(clk), .RN(n3023), .Q(
        \CACHE[4][37] ), .QN(n1198) );
  DFFRX1 \CACHE_reg[4][36]  ( .D(n2437), .CK(clk), .RN(n3038), .Q(
        \CACHE[4][36] ), .QN(n1197) );
  DFFRX1 \CACHE_reg[4][35]  ( .D(n2436), .CK(clk), .RN(n3026), .Q(
        \CACHE[4][35] ), .QN(n1196) );
  DFFRX1 \CACHE_reg[4][34]  ( .D(n2435), .CK(clk), .RN(n3028), .Q(
        \CACHE[4][34] ), .QN(n1195) );
  DFFRX1 \CACHE_reg[4][33]  ( .D(n2434), .CK(clk), .RN(n3038), .Q(
        \CACHE[4][33] ), .QN(n1194) );
  DFFRX1 \CACHE_reg[4][32]  ( .D(n2433), .CK(clk), .RN(n3031), .Q(
        \CACHE[4][32] ), .QN(n1193) );
  DFFRX1 \CACHE_reg[4][31]  ( .D(n2432), .CK(clk), .RN(n476), .Q(
        \CACHE[4][31] ), .QN(n1192) );
  DFFRX1 \CACHE_reg[4][30]  ( .D(n2431), .CK(clk), .RN(n478), .Q(
        \CACHE[4][30] ), .QN(n1191) );
  DFFRX1 \CACHE_reg[4][29]  ( .D(n2430), .CK(clk), .RN(n481), .Q(
        \CACHE[4][29] ), .QN(n1190) );
  DFFRX1 \CACHE_reg[4][28]  ( .D(n2429), .CK(clk), .RN(n484), .Q(
        \CACHE[4][28] ), .QN(n1189) );
  DFFRX1 \CACHE_reg[4][27]  ( .D(n2428), .CK(clk), .RN(n486), .Q(
        \CACHE[4][27] ), .QN(n1188) );
  DFFRX1 \CACHE_reg[4][26]  ( .D(n2427), .CK(clk), .RN(n489), .Q(
        \CACHE[4][26] ), .QN(n1187) );
  DFFRX1 \CACHE_reg[4][25]  ( .D(n2426), .CK(clk), .RN(n492), .Q(
        \CACHE[4][25] ), .QN(n1186) );
  DFFRX1 \CACHE_reg[4][24]  ( .D(n2425), .CK(clk), .RN(n494), .Q(
        \CACHE[4][24] ), .QN(n1185) );
  DFFRX1 \CACHE_reg[4][23]  ( .D(n2424), .CK(clk), .RN(n497), .Q(
        \CACHE[4][23] ), .QN(n1184) );
  DFFRX1 \CACHE_reg[4][22]  ( .D(n2423), .CK(clk), .RN(n500), .Q(
        \CACHE[4][22] ), .QN(n1183) );
  DFFRX1 \CACHE_reg[4][21]  ( .D(n2422), .CK(clk), .RN(n502), .Q(
        \CACHE[4][21] ), .QN(n1182) );
  DFFRX1 \CACHE_reg[4][20]  ( .D(n2421), .CK(clk), .RN(n505), .Q(
        \CACHE[4][20] ), .QN(n1181) );
  DFFRX1 \CACHE_reg[4][19]  ( .D(n2420), .CK(clk), .RN(n508), .Q(
        \CACHE[4][19] ), .QN(n1180) );
  DFFRX1 \CACHE_reg[4][18]  ( .D(n2419), .CK(clk), .RN(n3058), .Q(
        \CACHE[4][18] ), .QN(n1179) );
  DFFRX1 \CACHE_reg[4][17]  ( .D(n2418), .CK(clk), .RN(n510), .Q(
        \CACHE[4][17] ), .QN(n1178) );
  DFFRX1 \CACHE_reg[4][16]  ( .D(n2417), .CK(clk), .RN(n513), .Q(
        \CACHE[4][16] ), .QN(n1177) );
  DFFRX1 \CACHE_reg[4][15]  ( .D(n2416), .CK(clk), .RN(n516), .Q(
        \CACHE[4][15] ), .QN(n1176) );
  DFFRX1 \CACHE_reg[4][14]  ( .D(n2415), .CK(clk), .RN(n518), .Q(
        \CACHE[4][14] ), .QN(n1175) );
  DFFRX1 \CACHE_reg[4][13]  ( .D(n2414), .CK(clk), .RN(n521), .Q(
        \CACHE[4][13] ), .QN(n1174) );
  DFFRX1 \CACHE_reg[4][12]  ( .D(n2413), .CK(clk), .RN(n524), .Q(
        \CACHE[4][12] ), .QN(n1173) );
  DFFRX1 \CACHE_reg[4][11]  ( .D(n2412), .CK(clk), .RN(n526), .Q(
        \CACHE[4][11] ), .QN(n1172) );
  DFFRX1 \CACHE_reg[4][10]  ( .D(n2411), .CK(clk), .RN(n529), .Q(
        \CACHE[4][10] ), .QN(n1171) );
  DFFRX1 \CACHE_reg[4][9]  ( .D(n2410), .CK(clk), .RN(n532), .Q(\CACHE[4][9] ), 
        .QN(n1170) );
  DFFRX1 \CACHE_reg[4][8]  ( .D(n2409), .CK(clk), .RN(n534), .Q(\CACHE[4][8] ), 
        .QN(n1169) );
  DFFRX1 \CACHE_reg[4][7]  ( .D(n2408), .CK(clk), .RN(n537), .Q(\CACHE[4][7] ), 
        .QN(n1168) );
  DFFRX1 \CACHE_reg[4][6]  ( .D(n2407), .CK(clk), .RN(n540), .Q(\CACHE[4][6] ), 
        .QN(n1167) );
  DFFRX1 \CACHE_reg[4][5]  ( .D(n2406), .CK(clk), .RN(n3022), .Q(\CACHE[4][5] ), .QN(n1166) );
  DFFRX1 \CACHE_reg[4][4]  ( .D(n2405), .CK(clk), .RN(n3058), .Q(\CACHE[4][4] ), .QN(n1165) );
  DFFRX1 \CACHE_reg[4][3]  ( .D(n2404), .CK(clk), .RN(n3025), .Q(\CACHE[4][3] ), .QN(n1164) );
  DFFRX1 \CACHE_reg[4][2]  ( .D(n2403), .CK(clk), .RN(n3028), .Q(\CACHE[4][2] ), .QN(n1163) );
  DFFRX1 \CACHE_reg[4][1]  ( .D(n2402), .CK(clk), .RN(n3039), .Q(\CACHE[4][1] ), .QN(n1162) );
  DFFRX1 \CACHE_reg[4][0]  ( .D(n2401), .CK(clk), .RN(n3030), .Q(\CACHE[4][0] ), .QN(n1161) );
  DFFRX1 \CACHE_reg[0][154]  ( .D(n1935), .CK(clk), .RN(n3057), .Q(
        \CACHE[0][154] ), .QN(n695) );
  DFFRX1 \CACHE_reg[0][153]  ( .D(n1934), .CK(clk), .RN(n3057), .Q(
        \CACHE[0][153] ), .QN(n694) );
  DFFRX1 \CACHE_reg[0][152]  ( .D(n1933), .CK(clk), .RN(n3056), .Q(
        \CACHE[0][152] ), .QN(n693) );
  DFFRX1 \CACHE_reg[0][151]  ( .D(n1932), .CK(clk), .RN(n3040), .Q(
        \CACHE[0][151] ), .QN(n692) );
  DFFRX1 \CACHE_reg[0][150]  ( .D(n1931), .CK(clk), .RN(n3041), .Q(
        \CACHE[0][150] ), .QN(n691) );
  DFFRX1 \CACHE_reg[0][149]  ( .D(n1930), .CK(clk), .RN(n3041), .Q(
        \CACHE[0][149] ), .QN(n690) );
  DFFRX1 \CACHE_reg[0][148]  ( .D(n1929), .CK(clk), .RN(n3042), .Q(
        \CACHE[0][148] ), .QN(n689) );
  DFFRX1 \CACHE_reg[0][147]  ( .D(n1928), .CK(clk), .RN(n3043), .Q(
        \CACHE[0][147] ), .QN(n688) );
  DFFRX1 \CACHE_reg[0][146]  ( .D(n1927), .CK(clk), .RN(n3043), .Q(
        \CACHE[0][146] ), .QN(n687) );
  DFFRX1 \CACHE_reg[0][145]  ( .D(n1926), .CK(clk), .RN(n3044), .Q(
        \CACHE[0][145] ), .QN(n686) );
  DFFRX1 \CACHE_reg[0][144]  ( .D(n1925), .CK(clk), .RN(n3045), .Q(
        \CACHE[0][144] ), .QN(n685) );
  DFFRX1 \CACHE_reg[0][143]  ( .D(n1924), .CK(clk), .RN(n3045), .Q(
        \CACHE[0][143] ), .QN(n684) );
  DFFRX1 \CACHE_reg[0][142]  ( .D(n1923), .CK(clk), .RN(n3046), .Q(
        \CACHE[0][142] ), .QN(n683) );
  DFFRX1 \CACHE_reg[0][141]  ( .D(n1922), .CK(clk), .RN(n3047), .Q(
        \CACHE[0][141] ), .QN(n682) );
  DFFRX1 \CACHE_reg[0][140]  ( .D(n1921), .CK(clk), .RN(n3047), .Q(
        \CACHE[0][140] ), .QN(n681) );
  DFFRX1 \CACHE_reg[0][139]  ( .D(n1920), .CK(clk), .RN(n3048), .Q(
        \CACHE[0][139] ), .QN(n680) );
  DFFRX1 \CACHE_reg[0][138]  ( .D(n1919), .CK(clk), .RN(n3049), .Q(
        \CACHE[0][138] ), .QN(n679) );
  DFFRX1 \CACHE_reg[0][137]  ( .D(n1918), .CK(clk), .RN(n3049), .Q(
        \CACHE[0][137] ), .QN(n678) );
  DFFRX1 \CACHE_reg[0][136]  ( .D(n1917), .CK(clk), .RN(n3050), .Q(
        \CACHE[0][136] ), .QN(n677) );
  DFFRX1 \CACHE_reg[0][135]  ( .D(n1916), .CK(clk), .RN(n3051), .Q(
        \CACHE[0][135] ), .QN(n676) );
  DFFRX1 \CACHE_reg[0][134]  ( .D(n1915), .CK(clk), .RN(n3051), .Q(
        \CACHE[0][134] ), .QN(n675) );
  DFFRX1 \CACHE_reg[0][133]  ( .D(n1914), .CK(clk), .RN(n3052), .Q(
        \CACHE[0][133] ), .QN(n674) );
  DFFRX1 \CACHE_reg[0][132]  ( .D(n1913), .CK(clk), .RN(n3053), .Q(
        \CACHE[0][132] ), .QN(n673) );
  DFFRX1 \CACHE_reg[0][131]  ( .D(n1912), .CK(clk), .RN(n3053), .Q(
        \CACHE[0][131] ), .QN(n672) );
  DFFRX1 \CACHE_reg[0][130]  ( .D(n1911), .CK(clk), .RN(n3054), .Q(
        \CACHE[0][130] ), .QN(n671) );
  DFFRX1 \CACHE_reg[0][129]  ( .D(n1910), .CK(clk), .RN(n3055), .Q(
        \CACHE[0][129] ), .QN(n670) );
  DFFRX1 \CACHE_reg[0][128]  ( .D(n1909), .CK(clk), .RN(n3055), .Q(
        \CACHE[0][128] ), .QN(n669) );
  DFFRX1 \CACHE_reg[0][127]  ( .D(n1908), .CK(clk), .RN(n478), .Q(
        \CACHE[0][127] ), .QN(n668) );
  DFFRX1 \CACHE_reg[0][126]  ( .D(n1907), .CK(clk), .RN(n481), .Q(
        \CACHE[0][126] ), .QN(n667) );
  DFFRX1 \CACHE_reg[0][125]  ( .D(n1906), .CK(clk), .RN(n483), .Q(
        \CACHE[0][125] ), .QN(n666) );
  DFFRX1 \CACHE_reg[0][124]  ( .D(n1905), .CK(clk), .RN(n486), .Q(
        \CACHE[0][124] ), .QN(n665) );
  DFFRX1 \CACHE_reg[0][123]  ( .D(n1904), .CK(clk), .RN(n489), .Q(
        \CACHE[0][123] ), .QN(n664) );
  DFFRX1 \CACHE_reg[0][122]  ( .D(n1903), .CK(clk), .RN(n491), .Q(
        \CACHE[0][122] ), .QN(n663) );
  DFFRX1 \CACHE_reg[0][121]  ( .D(n1902), .CK(clk), .RN(n494), .Q(
        \CACHE[0][121] ), .QN(n662) );
  DFFRX1 \CACHE_reg[0][120]  ( .D(n1901), .CK(clk), .RN(n497), .Q(
        \CACHE[0][120] ), .QN(n661) );
  DFFRX1 \CACHE_reg[0][119]  ( .D(n1900), .CK(clk), .RN(n499), .Q(
        \CACHE[0][119] ), .QN(n660) );
  DFFRX1 \CACHE_reg[0][118]  ( .D(n1899), .CK(clk), .RN(n502), .Q(
        \CACHE[0][118] ), .QN(n659) );
  DFFRX1 \CACHE_reg[0][117]  ( .D(n1898), .CK(clk), .RN(n505), .Q(
        \CACHE[0][117] ), .QN(n658) );
  DFFRX1 \CACHE_reg[0][116]  ( .D(n1897), .CK(clk), .RN(n507), .Q(
        \CACHE[0][116] ), .QN(n657) );
  DFFRX1 \CACHE_reg[0][115]  ( .D(n1896), .CK(clk), .RN(n510), .Q(
        \CACHE[0][115] ), .QN(n656) );
  DFFRX1 \CACHE_reg[0][114]  ( .D(n1895), .CK(clk), .RN(n3033), .Q(
        \CACHE[0][114] ), .QN(n655) );
  DFFRX1 \CACHE_reg[0][113]  ( .D(n1894), .CK(clk), .RN(n513), .Q(
        \CACHE[0][113] ), .QN(n654) );
  DFFRX1 \CACHE_reg[0][112]  ( .D(n1893), .CK(clk), .RN(n515), .Q(
        \CACHE[0][112] ), .QN(n653) );
  DFFRX1 \CACHE_reg[0][111]  ( .D(n1892), .CK(clk), .RN(n518), .Q(
        \CACHE[0][111] ), .QN(n652) );
  DFFRX1 \CACHE_reg[0][110]  ( .D(n1891), .CK(clk), .RN(n521), .Q(
        \CACHE[0][110] ), .QN(n651) );
  DFFRX1 \CACHE_reg[0][109]  ( .D(n1890), .CK(clk), .RN(n523), .Q(
        \CACHE[0][109] ), .QN(n650) );
  DFFRX1 \CACHE_reg[0][108]  ( .D(n1889), .CK(clk), .RN(n526), .Q(
        \CACHE[0][108] ), .QN(n649) );
  DFFRX1 \CACHE_reg[0][107]  ( .D(n1888), .CK(clk), .RN(n529), .Q(
        \CACHE[0][107] ), .QN(n648) );
  DFFRX1 \CACHE_reg[0][106]  ( .D(n1887), .CK(clk), .RN(n531), .Q(
        \CACHE[0][106] ), .QN(n647) );
  DFFRX1 \CACHE_reg[0][105]  ( .D(n1886), .CK(clk), .RN(n534), .Q(
        \CACHE[0][105] ), .QN(n646) );
  DFFRX1 \CACHE_reg[0][104]  ( .D(n1885), .CK(clk), .RN(n537), .Q(
        \CACHE[0][104] ), .QN(n645) );
  DFFRX1 \CACHE_reg[0][103]  ( .D(n1884), .CK(clk), .RN(n539), .Q(
        \CACHE[0][103] ), .QN(n644) );
  DFFRX1 \CACHE_reg[0][102]  ( .D(n1883), .CK(clk), .RN(n3022), .Q(
        \CACHE[0][102] ), .QN(n643) );
  DFFRX1 \CACHE_reg[0][101]  ( .D(n1882), .CK(clk), .RN(n3025), .Q(
        \CACHE[0][101] ), .QN(n642) );
  DFFRX1 \CACHE_reg[0][100]  ( .D(n1881), .CK(clk), .RN(n3034), .Q(
        \CACHE[0][100] ), .QN(n641) );
  DFFRX1 \CACHE_reg[0][99]  ( .D(n1880), .CK(clk), .RN(n3027), .Q(
        \CACHE[0][99] ), .QN(n640) );
  DFFRX1 \CACHE_reg[0][98]  ( .D(n1879), .CK(clk), .RN(n3030), .Q(
        \CACHE[0][98] ), .QN(n639) );
  DFFRX1 \CACHE_reg[0][97]  ( .D(n1878), .CK(clk), .RN(n3035), .Q(
        \CACHE[0][97] ), .QN(n638) );
  DFFRX1 \CACHE_reg[0][96]  ( .D(n1877), .CK(clk), .RN(n3033), .Q(
        \CACHE[0][96] ), .QN(n637) );
  DFFRX1 \CACHE_reg[0][95]  ( .D(n1876), .CK(clk), .RN(n477), .Q(
        \CACHE[0][95] ), .QN(n636) );
  DFFRX1 \CACHE_reg[0][94]  ( .D(n1875), .CK(clk), .RN(n480), .Q(
        \CACHE[0][94] ), .QN(n635) );
  DFFRX1 \CACHE_reg[0][93]  ( .D(n1874), .CK(clk), .RN(n483), .Q(
        \CACHE[0][93] ), .QN(n634) );
  DFFRX1 \CACHE_reg[0][92]  ( .D(n1873), .CK(clk), .RN(n485), .Q(
        \CACHE[0][92] ), .QN(n633) );
  DFFRX1 \CACHE_reg[0][91]  ( .D(n1872), .CK(clk), .RN(n488), .Q(
        \CACHE[0][91] ), .QN(n632) );
  DFFRX1 \CACHE_reg[0][90]  ( .D(n1871), .CK(clk), .RN(n491), .Q(
        \CACHE[0][90] ), .QN(n631) );
  DFFRX1 \CACHE_reg[0][89]  ( .D(n1870), .CK(clk), .RN(n493), .Q(
        \CACHE[0][89] ), .QN(n630) );
  DFFRX1 \CACHE_reg[0][88]  ( .D(n1869), .CK(clk), .RN(n496), .Q(
        \CACHE[0][88] ), .QN(n629) );
  DFFRX1 \CACHE_reg[0][87]  ( .D(n1868), .CK(clk), .RN(n499), .Q(
        \CACHE[0][87] ), .QN(n628) );
  DFFRX1 \CACHE_reg[0][86]  ( .D(n1867), .CK(clk), .RN(n501), .Q(
        \CACHE[0][86] ), .QN(n627) );
  DFFRX1 \CACHE_reg[0][85]  ( .D(n1866), .CK(clk), .RN(n504), .Q(
        \CACHE[0][85] ), .QN(n626) );
  DFFRX1 \CACHE_reg[0][84]  ( .D(n1865), .CK(clk), .RN(n507), .Q(
        \CACHE[0][84] ), .QN(n625) );
  DFFRX1 \CACHE_reg[0][83]  ( .D(n1864), .CK(clk), .RN(n509), .Q(
        \CACHE[0][83] ), .QN(n624) );
  DFFRX1 \CACHE_reg[0][82]  ( .D(n1863), .CK(clk), .RN(n3035), .Q(
        \CACHE[0][82] ), .QN(n623) );
  DFFRX1 \CACHE_reg[0][81]  ( .D(n1862), .CK(clk), .RN(n512), .Q(
        \CACHE[0][81] ), .QN(n622) );
  DFFRX1 \CACHE_reg[0][80]  ( .D(n1861), .CK(clk), .RN(n515), .Q(
        \CACHE[0][80] ), .QN(n621) );
  DFFRX1 \CACHE_reg[0][79]  ( .D(n1860), .CK(clk), .RN(n517), .Q(
        \CACHE[0][79] ), .QN(n620) );
  DFFRX1 \CACHE_reg[0][78]  ( .D(n1859), .CK(clk), .RN(n520), .Q(
        \CACHE[0][78] ), .QN(n619) );
  DFFRX1 \CACHE_reg[0][77]  ( .D(n1858), .CK(clk), .RN(n523), .Q(
        \CACHE[0][77] ), .QN(n618) );
  DFFRX1 \CACHE_reg[0][76]  ( .D(n1857), .CK(clk), .RN(n525), .Q(
        \CACHE[0][76] ), .QN(n617) );
  DFFRX1 \CACHE_reg[0][75]  ( .D(n1856), .CK(clk), .RN(n528), .Q(
        \CACHE[0][75] ), .QN(n616) );
  DFFRX1 \CACHE_reg[0][74]  ( .D(n1855), .CK(clk), .RN(n531), .Q(
        \CACHE[0][74] ), .QN(n615) );
  DFFRX1 \CACHE_reg[0][73]  ( .D(n1854), .CK(clk), .RN(n533), .Q(
        \CACHE[0][73] ), .QN(n614) );
  DFFRX1 \CACHE_reg[0][72]  ( .D(n1853), .CK(clk), .RN(n536), .Q(
        \CACHE[0][72] ), .QN(n613) );
  DFFRX1 \CACHE_reg[0][71]  ( .D(n1852), .CK(clk), .RN(n539), .Q(
        \CACHE[0][71] ), .QN(n612) );
  DFFRX1 \CACHE_reg[0][70]  ( .D(n1851), .CK(clk), .RN(n3020), .Q(
        \CACHE[0][70] ), .QN(n611) );
  DFFRX1 \CACHE_reg[0][69]  ( .D(n1850), .CK(clk), .RN(n3024), .Q(
        \CACHE[0][69] ), .QN(n610) );
  DFFRX1 \CACHE_reg[0][68]  ( .D(n1849), .CK(clk), .RN(n3036), .Q(
        \CACHE[0][68] ), .QN(n609) );
  DFFRX1 \CACHE_reg[0][67]  ( .D(n1848), .CK(clk), .RN(n3027), .Q(
        \CACHE[0][67] ), .QN(n608) );
  DFFRX1 \CACHE_reg[0][66]  ( .D(n1847), .CK(clk), .RN(n3029), .Q(
        \CACHE[0][66] ), .QN(n607) );
  DFFRX1 \CACHE_reg[0][65]  ( .D(n1846), .CK(clk), .RN(n3037), .Q(
        \CACHE[0][65] ), .QN(n606) );
  DFFRX1 \CACHE_reg[0][64]  ( .D(n1845), .CK(clk), .RN(n3032), .Q(
        \CACHE[0][64] ), .QN(n605) );
  DFFRX1 \CACHE_reg[0][63]  ( .D(n1844), .CK(clk), .RN(n477), .Q(
        \CACHE[0][63] ), .QN(n604) );
  DFFRX1 \CACHE_reg[0][62]  ( .D(n1843), .CK(clk), .RN(n479), .Q(
        \CACHE[0][62] ), .QN(n603) );
  DFFRX1 \CACHE_reg[0][61]  ( .D(n1842), .CK(clk), .RN(n482), .Q(
        \CACHE[0][61] ), .QN(n602) );
  DFFRX1 \CACHE_reg[0][60]  ( .D(n1841), .CK(clk), .RN(n485), .Q(
        \CACHE[0][60] ), .QN(n601) );
  DFFRX1 \CACHE_reg[0][59]  ( .D(n1840), .CK(clk), .RN(n487), .Q(
        \CACHE[0][59] ), .QN(n600) );
  DFFRX1 \CACHE_reg[0][58]  ( .D(n1839), .CK(clk), .RN(n490), .Q(
        \CACHE[0][58] ), .QN(n599) );
  DFFRX1 \CACHE_reg[0][57]  ( .D(n1838), .CK(clk), .RN(n493), .Q(
        \CACHE[0][57] ), .QN(n598) );
  DFFRX1 \CACHE_reg[0][56]  ( .D(n1837), .CK(clk), .RN(n495), .Q(
        \CACHE[0][56] ), .QN(n597) );
  DFFRX1 \CACHE_reg[0][55]  ( .D(n1836), .CK(clk), .RN(n498), .Q(
        \CACHE[0][55] ), .QN(n596) );
  DFFRX1 \CACHE_reg[0][54]  ( .D(n1835), .CK(clk), .RN(n501), .Q(
        \CACHE[0][54] ), .QN(n595) );
  DFFRX1 \CACHE_reg[0][53]  ( .D(n1834), .CK(clk), .RN(n503), .Q(
        \CACHE[0][53] ), .QN(n594) );
  DFFRX1 \CACHE_reg[0][52]  ( .D(n1833), .CK(clk), .RN(n506), .Q(
        \CACHE[0][52] ), .QN(n593) );
  DFFRX1 \CACHE_reg[0][51]  ( .D(n1832), .CK(clk), .RN(n509), .Q(
        \CACHE[0][51] ), .QN(n592) );
  DFFRX1 \CACHE_reg[0][50]  ( .D(n1831), .CK(clk), .RN(n3037), .Q(
        \CACHE[0][50] ), .QN(n591) );
  DFFRX1 \CACHE_reg[0][49]  ( .D(n1830), .CK(clk), .RN(n511), .Q(
        \CACHE[0][49] ), .QN(n590) );
  DFFRX1 \CACHE_reg[0][48]  ( .D(n1829), .CK(clk), .RN(n514), .Q(
        \CACHE[0][48] ), .QN(n589) );
  DFFRX1 \CACHE_reg[0][47]  ( .D(n1828), .CK(clk), .RN(n517), .Q(
        \CACHE[0][47] ), .QN(n588) );
  DFFRX1 \CACHE_reg[0][46]  ( .D(n1827), .CK(clk), .RN(n519), .Q(
        \CACHE[0][46] ), .QN(n587) );
  DFFRX1 \CACHE_reg[0][45]  ( .D(n1826), .CK(clk), .RN(n522), .Q(
        \CACHE[0][45] ), .QN(n586) );
  DFFRX1 \CACHE_reg[0][44]  ( .D(n1825), .CK(clk), .RN(n525), .Q(
        \CACHE[0][44] ), .QN(n585) );
  DFFRX1 \CACHE_reg[0][43]  ( .D(n1824), .CK(clk), .RN(n527), .Q(
        \CACHE[0][43] ), .QN(n584) );
  DFFRX1 \CACHE_reg[0][42]  ( .D(n1823), .CK(clk), .RN(n530), .Q(
        \CACHE[0][42] ), .QN(n583) );
  DFFRX1 \CACHE_reg[0][41]  ( .D(n1822), .CK(clk), .RN(n533), .Q(
        \CACHE[0][41] ), .QN(n582) );
  DFFRX1 \CACHE_reg[0][40]  ( .D(n1821), .CK(clk), .RN(n535), .Q(
        \CACHE[0][40] ), .QN(n581) );
  DFFRX1 \CACHE_reg[0][39]  ( .D(n1820), .CK(clk), .RN(n538), .Q(
        \CACHE[0][39] ), .QN(n580) );
  DFFRX1 \CACHE_reg[0][38]  ( .D(n1819), .CK(clk), .RN(n3020), .Q(
        \CACHE[0][38] ), .QN(n579) );
  DFFRX1 \CACHE_reg[0][37]  ( .D(n1818), .CK(clk), .RN(n3023), .Q(
        \CACHE[0][37] ), .QN(n578) );
  DFFRX1 \CACHE_reg[0][36]  ( .D(n1817), .CK(clk), .RN(n3038), .Q(
        \CACHE[0][36] ), .QN(n577) );
  DFFRX1 \CACHE_reg[0][35]  ( .D(n1816), .CK(clk), .RN(n3026), .Q(
        \CACHE[0][35] ), .QN(n576) );
  DFFRX1 \CACHE_reg[0][34]  ( .D(n1815), .CK(clk), .RN(n3029), .Q(
        \CACHE[0][34] ), .QN(n575) );
  DFFRX1 \CACHE_reg[0][33]  ( .D(n1814), .CK(clk), .RN(n3039), .Q(
        \CACHE[0][33] ), .QN(n574) );
  DFFRX1 \CACHE_reg[0][32]  ( .D(n1813), .CK(clk), .RN(n3031), .Q(
        \CACHE[0][32] ), .QN(n573) );
  DFFRX1 \CACHE_reg[0][31]  ( .D(n1812), .CK(clk), .RN(n476), .Q(
        \CACHE[0][31] ), .QN(n572) );
  DFFRX1 \CACHE_reg[0][30]  ( .D(n1811), .CK(clk), .RN(n479), .Q(
        \CACHE[0][30] ), .QN(n571) );
  DFFRX1 \CACHE_reg[0][29]  ( .D(n1810), .CK(clk), .RN(n481), .Q(
        \CACHE[0][29] ), .QN(n570) );
  DFFRX1 \CACHE_reg[0][28]  ( .D(n1809), .CK(clk), .RN(n484), .Q(
        \CACHE[0][28] ), .QN(n569) );
  DFFRX1 \CACHE_reg[0][27]  ( .D(n1808), .CK(clk), .RN(n487), .Q(
        \CACHE[0][27] ), .QN(n568) );
  DFFRX1 \CACHE_reg[0][26]  ( .D(n1807), .CK(clk), .RN(n489), .Q(
        \CACHE[0][26] ), .QN(n567) );
  DFFRX1 \CACHE_reg[0][25]  ( .D(n1806), .CK(clk), .RN(n492), .Q(
        \CACHE[0][25] ), .QN(n566) );
  DFFRX1 \CACHE_reg[0][24]  ( .D(n1805), .CK(clk), .RN(n495), .Q(
        \CACHE[0][24] ), .QN(n565) );
  DFFRX1 \CACHE_reg[0][23]  ( .D(n1804), .CK(clk), .RN(n497), .Q(
        \CACHE[0][23] ), .QN(n564) );
  DFFRX1 \CACHE_reg[0][22]  ( .D(n1803), .CK(clk), .RN(n500), .Q(
        \CACHE[0][22] ), .QN(n563) );
  DFFRX1 \CACHE_reg[0][21]  ( .D(n1802), .CK(clk), .RN(n503), .Q(
        \CACHE[0][21] ), .QN(n562) );
  DFFRX1 \CACHE_reg[0][20]  ( .D(n1801), .CK(clk), .RN(n505), .Q(
        \CACHE[0][20] ), .QN(n561) );
  DFFRX1 \CACHE_reg[0][19]  ( .D(n1800), .CK(clk), .RN(n508), .Q(
        \CACHE[0][19] ), .QN(n560) );
  DFFRX1 \CACHE_reg[0][18]  ( .D(n1799), .CK(clk), .RN(n3059), .Q(
        \CACHE[0][18] ), .QN(n559) );
  DFFRX1 \CACHE_reg[0][17]  ( .D(n1798), .CK(clk), .RN(n511), .Q(
        \CACHE[0][17] ), .QN(n558) );
  DFFRX1 \CACHE_reg[0][16]  ( .D(n1797), .CK(clk), .RN(n513), .Q(
        \CACHE[0][16] ), .QN(n557) );
  DFFRX1 \CACHE_reg[0][15]  ( .D(n1796), .CK(clk), .RN(n516), .Q(
        \CACHE[0][15] ), .QN(n556) );
  DFFRX1 \CACHE_reg[0][14]  ( .D(n1795), .CK(clk), .RN(n519), .Q(
        \CACHE[0][14] ), .QN(n555) );
  DFFRX1 \CACHE_reg[0][13]  ( .D(n1794), .CK(clk), .RN(n521), .Q(
        \CACHE[0][13] ), .QN(n554) );
  DFFRX1 \CACHE_reg[0][12]  ( .D(n1793), .CK(clk), .RN(n524), .Q(
        \CACHE[0][12] ), .QN(n553) );
  DFFRX1 \CACHE_reg[0][11]  ( .D(n1792), .CK(clk), .RN(n527), .Q(
        \CACHE[0][11] ), .QN(n552) );
  DFFRX1 \CACHE_reg[0][10]  ( .D(n1791), .CK(clk), .RN(n529), .Q(
        \CACHE[0][10] ), .QN(n551) );
  DFFRX1 \CACHE_reg[0][9]  ( .D(n1790), .CK(clk), .RN(n532), .Q(\CACHE[0][9] ), 
        .QN(n550) );
  DFFRX1 \CACHE_reg[0][8]  ( .D(n1789), .CK(clk), .RN(n535), .Q(\CACHE[0][8] ), 
        .QN(n549) );
  DFFRX1 \CACHE_reg[0][7]  ( .D(n1788), .CK(clk), .RN(n537), .Q(\CACHE[0][7] ), 
        .QN(n548) );
  DFFRX1 \CACHE_reg[0][6]  ( .D(n1787), .CK(clk), .RN(n540), .Q(\CACHE[0][6] ), 
        .QN(n547) );
  DFFRX1 \CACHE_reg[0][5]  ( .D(n1786), .CK(clk), .RN(n3023), .Q(\CACHE[0][5] ), .QN(n546) );
  DFFRX1 \CACHE_reg[0][4]  ( .D(n1785), .CK(clk), .RN(n3058), .Q(\CACHE[0][4] ), .QN(n545) );
  DFFRX1 \CACHE_reg[0][3]  ( .D(n1784), .CK(clk), .RN(n3025), .Q(\CACHE[0][3] ), .QN(n544) );
  DFFRX1 \CACHE_reg[0][2]  ( .D(n1783), .CK(clk), .RN(n3028), .Q(\CACHE[0][2] ), .QN(n543) );
  DFFRX1 \CACHE_reg[0][1]  ( .D(n1782), .CK(clk), .RN(n3039), .Q(\CACHE[0][1] ), .QN(n542) );
  DFFRX1 \CACHE_reg[0][0]  ( .D(n1781), .CK(clk), .RN(n3031), .Q(\CACHE[0][0] ), .QN(n541) );
  DFFRX1 \CACHE_reg[6][154]  ( .D(n2865), .CK(clk), .RN(n3057), .Q(
        \CACHE[6][154] ), .QN(n1625) );
  DFFRX1 \CACHE_reg[6][153]  ( .D(n2864), .CK(clk), .RN(n3056), .Q(
        \CACHE[6][153] ), .QN(n1624) );
  DFFRX1 \CACHE_reg[6][152]  ( .D(n2863), .CK(clk), .RN(n3056), .Q(
        \CACHE[6][152] ), .QN(n1623) );
  DFFRX1 \CACHE_reg[6][151]  ( .D(n2862), .CK(clk), .RN(n3040), .Q(
        \CACHE[6][151] ), .QN(n1622) );
  DFFRX1 \CACHE_reg[6][150]  ( .D(n2861), .CK(clk), .RN(n3040), .Q(
        \CACHE[6][150] ), .QN(n1621) );
  DFFRX1 \CACHE_reg[6][149]  ( .D(n2860), .CK(clk), .RN(n3041), .Q(
        \CACHE[6][149] ), .QN(n1620) );
  DFFRX1 \CACHE_reg[6][148]  ( .D(n2859), .CK(clk), .RN(n3042), .Q(
        \CACHE[6][148] ), .QN(n1619) );
  DFFRX1 \CACHE_reg[6][147]  ( .D(n2858), .CK(clk), .RN(n3042), .Q(
        \CACHE[6][147] ), .QN(n1618) );
  DFFRX1 \CACHE_reg[6][146]  ( .D(n2857), .CK(clk), .RN(n3043), .Q(
        \CACHE[6][146] ), .QN(n1617) );
  DFFRX1 \CACHE_reg[6][145]  ( .D(n2856), .CK(clk), .RN(n3044), .Q(
        \CACHE[6][145] ), .QN(n1616) );
  DFFRX1 \CACHE_reg[6][144]  ( .D(n2855), .CK(clk), .RN(n3044), .Q(
        \CACHE[6][144] ), .QN(n1615) );
  DFFRX1 \CACHE_reg[6][143]  ( .D(n2854), .CK(clk), .RN(n3045), .Q(
        \CACHE[6][143] ), .QN(n1614) );
  DFFRX1 \CACHE_reg[6][142]  ( .D(n2853), .CK(clk), .RN(n3046), .Q(
        \CACHE[6][142] ), .QN(n1613) );
  DFFRX1 \CACHE_reg[6][141]  ( .D(n2852), .CK(clk), .RN(n3046), .Q(
        \CACHE[6][141] ), .QN(n1612) );
  DFFRX1 \CACHE_reg[6][140]  ( .D(n2851), .CK(clk), .RN(n3047), .Q(
        \CACHE[6][140] ), .QN(n1611) );
  DFFRX1 \CACHE_reg[6][139]  ( .D(n2850), .CK(clk), .RN(n3048), .Q(
        \CACHE[6][139] ), .QN(n1610) );
  DFFRX1 \CACHE_reg[6][138]  ( .D(n2849), .CK(clk), .RN(n3048), .Q(
        \CACHE[6][138] ), .QN(n1609) );
  DFFRX1 \CACHE_reg[6][137]  ( .D(n2848), .CK(clk), .RN(n3049), .Q(
        \CACHE[6][137] ), .QN(n1608) );
  DFFRX1 \CACHE_reg[6][136]  ( .D(n2847), .CK(clk), .RN(n3050), .Q(
        \CACHE[6][136] ), .QN(n1607) );
  DFFRX1 \CACHE_reg[6][135]  ( .D(n2846), .CK(clk), .RN(n3050), .Q(
        \CACHE[6][135] ), .QN(n1606) );
  DFFRX1 \CACHE_reg[6][134]  ( .D(n2845), .CK(clk), .RN(n3051), .Q(
        \CACHE[6][134] ), .QN(n1605) );
  DFFRX1 \CACHE_reg[6][133]  ( .D(n2844), .CK(clk), .RN(n3052), .Q(
        \CACHE[6][133] ), .QN(n1604) );
  DFFRX1 \CACHE_reg[6][132]  ( .D(n2843), .CK(clk), .RN(n3052), .Q(
        \CACHE[6][132] ), .QN(n1603) );
  DFFRX1 \CACHE_reg[6][131]  ( .D(n2842), .CK(clk), .RN(n3053), .Q(
        \CACHE[6][131] ), .QN(n1602) );
  DFFRX1 \CACHE_reg[6][130]  ( .D(n2841), .CK(clk), .RN(n3054), .Q(
        \CACHE[6][130] ), .QN(n1601) );
  DFFRX1 \CACHE_reg[6][129]  ( .D(n2840), .CK(clk), .RN(n3054), .Q(
        \CACHE[6][129] ), .QN(n1600) );
  DFFRX1 \CACHE_reg[6][128]  ( .D(n2839), .CK(clk), .RN(n3055), .Q(
        \CACHE[6][128] ), .QN(n1599) );
  DFFRX1 \CACHE_reg[6][127]  ( .D(n2838), .CK(clk), .RN(n478), .Q(
        \CACHE[6][127] ), .QN(n1598) );
  DFFRX1 \CACHE_reg[6][126]  ( .D(n2837), .CK(clk), .RN(n480), .Q(
        \CACHE[6][126] ), .QN(n1597) );
  DFFRX1 \CACHE_reg[6][125]  ( .D(n2836), .CK(clk), .RN(n483), .Q(
        \CACHE[6][125] ), .QN(n1596) );
  DFFRX1 \CACHE_reg[6][124]  ( .D(n2835), .CK(clk), .RN(n486), .Q(
        \CACHE[6][124] ), .QN(n1595) );
  DFFRX1 \CACHE_reg[6][123]  ( .D(n2834), .CK(clk), .RN(n488), .Q(
        \CACHE[6][123] ), .QN(n1594) );
  DFFRX1 \CACHE_reg[6][122]  ( .D(n2833), .CK(clk), .RN(n491), .Q(
        \CACHE[6][122] ), .QN(n1593) );
  DFFRX1 \CACHE_reg[6][121]  ( .D(n2832), .CK(clk), .RN(n494), .Q(
        \CACHE[6][121] ), .QN(n1592) );
  DFFRX1 \CACHE_reg[6][120]  ( .D(n2831), .CK(clk), .RN(n496), .Q(
        \CACHE[6][120] ), .QN(n1591) );
  DFFRX1 \CACHE_reg[6][119]  ( .D(n2830), .CK(clk), .RN(n499), .Q(
        \CACHE[6][119] ), .QN(n1590) );
  DFFRX1 \CACHE_reg[6][118]  ( .D(n2829), .CK(clk), .RN(n502), .Q(
        \CACHE[6][118] ), .QN(n1589) );
  DFFRX1 \CACHE_reg[6][117]  ( .D(n2828), .CK(clk), .RN(n504), .Q(
        \CACHE[6][117] ), .QN(n1588) );
  DFFRX1 \CACHE_reg[6][116]  ( .D(n2827), .CK(clk), .RN(n507), .Q(
        \CACHE[6][116] ), .QN(n1587) );
  DFFRX1 \CACHE_reg[6][115]  ( .D(n2826), .CK(clk), .RN(n510), .Q(
        \CACHE[6][115] ), .QN(n1586) );
  DFFRX1 \CACHE_reg[6][114]  ( .D(n2825), .CK(clk), .RN(n3033), .Q(
        \CACHE[6][114] ), .QN(n1585) );
  DFFRX1 \CACHE_reg[6][113]  ( .D(n2824), .CK(clk), .RN(n512), .Q(
        \CACHE[6][113] ), .QN(n1584) );
  DFFRX1 \CACHE_reg[6][112]  ( .D(n2823), .CK(clk), .RN(n515), .Q(
        \CACHE[6][112] ), .QN(n1583) );
  DFFRX1 \CACHE_reg[6][111]  ( .D(n2822), .CK(clk), .RN(n518), .Q(
        \CACHE[6][111] ), .QN(n1582) );
  DFFRX1 \CACHE_reg[6][110]  ( .D(n2821), .CK(clk), .RN(n520), .Q(
        \CACHE[6][110] ), .QN(n1581) );
  DFFRX1 \CACHE_reg[6][109]  ( .D(n2820), .CK(clk), .RN(n523), .Q(
        \CACHE[6][109] ), .QN(n1580) );
  DFFRX1 \CACHE_reg[6][108]  ( .D(n2819), .CK(clk), .RN(n526), .Q(
        \CACHE[6][108] ), .QN(n1579) );
  DFFRX1 \CACHE_reg[6][107]  ( .D(n2818), .CK(clk), .RN(n528), .Q(
        \CACHE[6][107] ), .QN(n1578) );
  DFFRX1 \CACHE_reg[6][106]  ( .D(n2817), .CK(clk), .RN(n531), .Q(
        \CACHE[6][106] ), .QN(n1577) );
  DFFRX1 \CACHE_reg[6][105]  ( .D(n2816), .CK(clk), .RN(n534), .Q(
        \CACHE[6][105] ), .QN(n1576) );
  DFFRX1 \CACHE_reg[6][104]  ( .D(n2815), .CK(clk), .RN(n536), .Q(
        \CACHE[6][104] ), .QN(n1575) );
  DFFRX1 \CACHE_reg[6][103]  ( .D(n2814), .CK(clk), .RN(n539), .Q(
        \CACHE[6][103] ), .QN(n1574) );
  DFFRX1 \CACHE_reg[6][102]  ( .D(n2813), .CK(clk), .RN(n3022), .Q(
        \CACHE[6][102] ), .QN(n1573) );
  DFFRX1 \CACHE_reg[6][101]  ( .D(n2812), .CK(clk), .RN(n3024), .Q(
        \CACHE[6][101] ), .QN(n1572) );
  DFFRX1 \CACHE_reg[6][100]  ( .D(n2811), .CK(clk), .RN(n3034), .Q(
        \CACHE[6][100] ), .QN(n1571) );
  DFFRX1 \CACHE_reg[6][99]  ( .D(n2810), .CK(clk), .RN(n3027), .Q(
        \CACHE[6][99] ), .QN(n1570) );
  DFFRX1 \CACHE_reg[6][98]  ( .D(n2809), .CK(clk), .RN(n3030), .Q(
        \CACHE[6][98] ), .QN(n1569) );
  DFFRX1 \CACHE_reg[6][97]  ( .D(n2808), .CK(clk), .RN(n3034), .Q(
        \CACHE[6][97] ), .QN(n1568) );
  DFFRX1 \CACHE_reg[6][96]  ( .D(n2807), .CK(clk), .RN(n3032), .Q(
        \CACHE[6][96] ), .QN(n1567) );
  DFFRX1 \CACHE_reg[6][95]  ( .D(n2806), .CK(clk), .RN(n477), .Q(
        \CACHE[6][95] ), .QN(n1566) );
  DFFRX1 \CACHE_reg[6][94]  ( .D(n2805), .CK(clk), .RN(n480), .Q(
        \CACHE[6][94] ), .QN(n1565) );
  DFFRX1 \CACHE_reg[6][93]  ( .D(n2804), .CK(clk), .RN(n482), .Q(
        \CACHE[6][93] ), .QN(n1564) );
  DFFRX1 \CACHE_reg[6][92]  ( .D(n2803), .CK(clk), .RN(n485), .Q(
        \CACHE[6][92] ), .QN(n1563) );
  DFFRX1 \CACHE_reg[6][91]  ( .D(n2802), .CK(clk), .RN(n488), .Q(
        \CACHE[6][91] ), .QN(n1562) );
  DFFRX1 \CACHE_reg[6][90]  ( .D(n2801), .CK(clk), .RN(n490), .Q(
        \CACHE[6][90] ), .QN(n1561) );
  DFFRX1 \CACHE_reg[6][89]  ( .D(n2800), .CK(clk), .RN(n493), .Q(
        \CACHE[6][89] ), .QN(n1560) );
  DFFRX1 \CACHE_reg[6][88]  ( .D(n2799), .CK(clk), .RN(n496), .Q(
        \CACHE[6][88] ), .QN(n1559) );
  DFFRX1 \CACHE_reg[6][87]  ( .D(n2798), .CK(clk), .RN(n498), .Q(
        \CACHE[6][87] ), .QN(n1558) );
  DFFRX1 \CACHE_reg[6][86]  ( .D(n2797), .CK(clk), .RN(n501), .Q(
        \CACHE[6][86] ), .QN(n1557) );
  DFFRX1 \CACHE_reg[6][85]  ( .D(n2796), .CK(clk), .RN(n504), .Q(
        \CACHE[6][85] ), .QN(n1556) );
  DFFRX1 \CACHE_reg[6][84]  ( .D(n2795), .CK(clk), .RN(n506), .Q(
        \CACHE[6][84] ), .QN(n1555) );
  DFFRX1 \CACHE_reg[6][83]  ( .D(n2794), .CK(clk), .RN(n509), .Q(
        \CACHE[6][83] ), .QN(n1554) );
  DFFRX1 \CACHE_reg[6][82]  ( .D(n2793), .CK(clk), .RN(n3035), .Q(
        \CACHE[6][82] ), .QN(n1553) );
  DFFRX1 \CACHE_reg[6][81]  ( .D(n2792), .CK(clk), .RN(n512), .Q(
        \CACHE[6][81] ), .QN(n1552) );
  DFFRX1 \CACHE_reg[6][80]  ( .D(n2791), .CK(clk), .RN(n514), .Q(
        \CACHE[6][80] ), .QN(n1551) );
  DFFRX1 \CACHE_reg[6][79]  ( .D(n2790), .CK(clk), .RN(n517), .Q(
        \CACHE[6][79] ), .QN(n1550) );
  DFFRX1 \CACHE_reg[6][78]  ( .D(n2789), .CK(clk), .RN(n520), .Q(
        \CACHE[6][78] ), .QN(n1549) );
  DFFRX1 \CACHE_reg[6][77]  ( .D(n2788), .CK(clk), .RN(n522), .Q(
        \CACHE[6][77] ), .QN(n1548) );
  DFFRX1 \CACHE_reg[6][76]  ( .D(n2787), .CK(clk), .RN(n525), .Q(
        \CACHE[6][76] ), .QN(n1547) );
  DFFRX1 \CACHE_reg[6][75]  ( .D(n2786), .CK(clk), .RN(n528), .Q(
        \CACHE[6][75] ), .QN(n1546) );
  DFFRX1 \CACHE_reg[6][74]  ( .D(n2785), .CK(clk), .RN(n530), .Q(
        \CACHE[6][74] ), .QN(n1545) );
  DFFRX1 \CACHE_reg[6][73]  ( .D(n2784), .CK(clk), .RN(n533), .Q(
        \CACHE[6][73] ), .QN(n1544) );
  DFFRX1 \CACHE_reg[6][72]  ( .D(n2783), .CK(clk), .RN(n536), .Q(
        \CACHE[6][72] ), .QN(n1543) );
  DFFRX1 \CACHE_reg[6][71]  ( .D(n2782), .CK(clk), .RN(n538), .Q(
        \CACHE[6][71] ), .QN(n1542) );
  DFFRX1 \CACHE_reg[6][70]  ( .D(n2781), .CK(clk), .RN(n3020), .Q(
        \CACHE[6][70] ), .QN(n1541) );
  DFFRX1 \CACHE_reg[6][69]  ( .D(n2780), .CK(clk), .RN(n3024), .Q(
        \CACHE[6][69] ), .QN(n1540) );
  DFFRX1 \CACHE_reg[6][68]  ( .D(n2779), .CK(clk), .RN(n3036), .Q(
        \CACHE[6][68] ), .QN(n1539) );
  DFFRX1 \CACHE_reg[6][67]  ( .D(n2778), .CK(clk), .RN(n3026), .Q(
        \CACHE[6][67] ), .QN(n1538) );
  DFFRX1 \CACHE_reg[6][66]  ( .D(n2777), .CK(clk), .RN(n3029), .Q(
        \CACHE[6][66] ), .QN(n1537) );
  DFFRX1 \CACHE_reg[6][65]  ( .D(n2776), .CK(clk), .RN(n3036), .Q(
        \CACHE[6][65] ), .QN(n1536) );
  DFFRX1 \CACHE_reg[6][64]  ( .D(n2775), .CK(clk), .RN(n3032), .Q(
        \CACHE[6][64] ), .QN(n1535) );
  DFFRX1 \CACHE_reg[6][63]  ( .D(n2774), .CK(clk), .RN(n476), .Q(
        \CACHE[6][63] ), .QN(n1534) );
  DFFRX1 \CACHE_reg[6][62]  ( .D(n2773), .CK(clk), .RN(n479), .Q(
        \CACHE[6][62] ), .QN(n1533) );
  DFFRX1 \CACHE_reg[6][61]  ( .D(n2772), .CK(clk), .RN(n482), .Q(
        \CACHE[6][61] ), .QN(n1532) );
  DFFRX1 \CACHE_reg[6][60]  ( .D(n2771), .CK(clk), .RN(n484), .Q(
        \CACHE[6][60] ), .QN(n1531) );
  DFFRX1 \CACHE_reg[6][59]  ( .D(n2770), .CK(clk), .RN(n487), .Q(
        \CACHE[6][59] ), .QN(n1530) );
  DFFRX1 \CACHE_reg[6][58]  ( .D(n2769), .CK(clk), .RN(n490), .Q(
        \CACHE[6][58] ), .QN(n1529) );
  DFFRX1 \CACHE_reg[6][57]  ( .D(n2768), .CK(clk), .RN(n492), .Q(
        \CACHE[6][57] ), .QN(n1528) );
  DFFRX1 \CACHE_reg[6][56]  ( .D(n2767), .CK(clk), .RN(n495), .Q(
        \CACHE[6][56] ), .QN(n1527) );
  DFFRX1 \CACHE_reg[6][55]  ( .D(n2766), .CK(clk), .RN(n498), .Q(
        \CACHE[6][55] ), .QN(n1526) );
  DFFRX1 \CACHE_reg[6][54]  ( .D(n2765), .CK(clk), .RN(n500), .Q(
        \CACHE[6][54] ), .QN(n1525) );
  DFFRX1 \CACHE_reg[6][53]  ( .D(n2764), .CK(clk), .RN(n503), .Q(
        \CACHE[6][53] ), .QN(n1524) );
  DFFRX1 \CACHE_reg[6][52]  ( .D(n2763), .CK(clk), .RN(n506), .Q(
        \CACHE[6][52] ), .QN(n1523) );
  DFFRX1 \CACHE_reg[6][51]  ( .D(n2762), .CK(clk), .RN(n508), .Q(
        \CACHE[6][51] ), .QN(n1522) );
  DFFRX1 \CACHE_reg[6][50]  ( .D(n2761), .CK(clk), .RN(n3037), .Q(
        \CACHE[6][50] ), .QN(n1521) );
  DFFRX1 \CACHE_reg[6][49]  ( .D(n2760), .CK(clk), .RN(n511), .Q(
        \CACHE[6][49] ), .QN(n1520) );
  DFFRX1 \CACHE_reg[6][48]  ( .D(n2759), .CK(clk), .RN(n514), .Q(
        \CACHE[6][48] ), .QN(n1519) );
  DFFRX1 \CACHE_reg[6][47]  ( .D(n2758), .CK(clk), .RN(n516), .Q(
        \CACHE[6][47] ), .QN(n1518) );
  DFFRX1 \CACHE_reg[6][46]  ( .D(n2757), .CK(clk), .RN(n519), .Q(
        \CACHE[6][46] ), .QN(n1517) );
  DFFRX1 \CACHE_reg[6][45]  ( .D(n2756), .CK(clk), .RN(n522), .Q(
        \CACHE[6][45] ), .QN(n1516) );
  DFFRX1 \CACHE_reg[6][44]  ( .D(n2755), .CK(clk), .RN(n524), .Q(
        \CACHE[6][44] ), .QN(n1515) );
  DFFRX1 \CACHE_reg[6][43]  ( .D(n2754), .CK(clk), .RN(n527), .Q(
        \CACHE[6][43] ), .QN(n1514) );
  DFFRX1 \CACHE_reg[6][42]  ( .D(n2753), .CK(clk), .RN(n530), .Q(
        \CACHE[6][42] ), .QN(n1513) );
  DFFRX1 \CACHE_reg[6][41]  ( .D(n2752), .CK(clk), .RN(n532), .Q(
        \CACHE[6][41] ), .QN(n1512) );
  DFFRX1 \CACHE_reg[6][40]  ( .D(n2751), .CK(clk), .RN(n535), .Q(
        \CACHE[6][40] ), .QN(n1511) );
  DFFRX1 \CACHE_reg[6][39]  ( .D(n2750), .CK(clk), .RN(n538), .Q(
        \CACHE[6][39] ), .QN(n1510) );
  DFFRX1 \CACHE_reg[6][38]  ( .D(n2749), .CK(clk), .RN(n540), .Q(
        \CACHE[6][38] ), .QN(n1509) );
  DFFRX1 \CACHE_reg[6][37]  ( .D(n2748), .CK(clk), .RN(n3023), .Q(
        \CACHE[6][37] ), .QN(n1508) );
  DFFRX1 \CACHE_reg[6][36]  ( .D(n2747), .CK(clk), .RN(n3038), .Q(
        \CACHE[6][36] ), .QN(n1507) );
  DFFRX1 \CACHE_reg[6][35]  ( .D(n2746), .CK(clk), .RN(n3026), .Q(
        \CACHE[6][35] ), .QN(n1506) );
  DFFRX1 \CACHE_reg[6][34]  ( .D(n2745), .CK(clk), .RN(n3028), .Q(
        \CACHE[6][34] ), .QN(n1505) );
  DFFRX1 \CACHE_reg[6][33]  ( .D(n2744), .CK(clk), .RN(n3038), .Q(
        \CACHE[6][33] ), .QN(n1504) );
  DFFRX1 \CACHE_reg[6][32]  ( .D(n2743), .CK(clk), .RN(n3031), .Q(
        \CACHE[6][32] ), .QN(n1503) );
  DFFRX1 \CACHE_reg[6][31]  ( .D(n2742), .CK(clk), .RN(n476), .Q(
        \CACHE[6][31] ), .QN(n1502) );
  DFFRX1 \CACHE_reg[6][30]  ( .D(n2741), .CK(clk), .RN(n478), .Q(
        \CACHE[6][30] ), .QN(n1501) );
  DFFRX1 \CACHE_reg[6][29]  ( .D(n2740), .CK(clk), .RN(n481), .Q(
        \CACHE[6][29] ), .QN(n1500) );
  DFFRX1 \CACHE_reg[6][28]  ( .D(n2739), .CK(clk), .RN(n484), .Q(
        \CACHE[6][28] ), .QN(n1499) );
  DFFRX1 \CACHE_reg[6][27]  ( .D(n2738), .CK(clk), .RN(n486), .Q(
        \CACHE[6][27] ), .QN(n1498) );
  DFFRX1 \CACHE_reg[6][26]  ( .D(n2737), .CK(clk), .RN(n489), .Q(
        \CACHE[6][26] ), .QN(n1497) );
  DFFRX1 \CACHE_reg[6][25]  ( .D(n2736), .CK(clk), .RN(n492), .Q(
        \CACHE[6][25] ), .QN(n1496) );
  DFFRX1 \CACHE_reg[6][24]  ( .D(n2735), .CK(clk), .RN(n494), .Q(
        \CACHE[6][24] ), .QN(n1495) );
  DFFRX1 \CACHE_reg[6][23]  ( .D(n2734), .CK(clk), .RN(n497), .Q(
        \CACHE[6][23] ), .QN(n1494) );
  DFFRX1 \CACHE_reg[6][22]  ( .D(n2733), .CK(clk), .RN(n500), .Q(
        \CACHE[6][22] ), .QN(n1493) );
  DFFRX1 \CACHE_reg[6][21]  ( .D(n2732), .CK(clk), .RN(n502), .Q(
        \CACHE[6][21] ), .QN(n1492) );
  DFFRX1 \CACHE_reg[6][20]  ( .D(n2731), .CK(clk), .RN(n505), .Q(
        \CACHE[6][20] ), .QN(n1491) );
  DFFRX1 \CACHE_reg[6][19]  ( .D(n2730), .CK(clk), .RN(n508), .Q(
        \CACHE[6][19] ), .QN(n1490) );
  DFFRX1 \CACHE_reg[6][18]  ( .D(n2729), .CK(clk), .RN(n3058), .Q(
        \CACHE[6][18] ), .QN(n1489) );
  DFFRX1 \CACHE_reg[6][17]  ( .D(n2728), .CK(clk), .RN(n510), .Q(
        \CACHE[6][17] ), .QN(n1488) );
  DFFRX1 \CACHE_reg[6][16]  ( .D(n2727), .CK(clk), .RN(n513), .Q(
        \CACHE[6][16] ), .QN(n1487) );
  DFFRX1 \CACHE_reg[6][15]  ( .D(n2726), .CK(clk), .RN(n516), .Q(
        \CACHE[6][15] ), .QN(n1486) );
  DFFRX1 \CACHE_reg[6][14]  ( .D(n2725), .CK(clk), .RN(n518), .Q(
        \CACHE[6][14] ), .QN(n1485) );
  DFFRX1 \CACHE_reg[6][13]  ( .D(n2724), .CK(clk), .RN(n521), .Q(
        \CACHE[6][13] ), .QN(n1484) );
  DFFRX1 \CACHE_reg[6][12]  ( .D(n2723), .CK(clk), .RN(n524), .Q(
        \CACHE[6][12] ), .QN(n1483) );
  DFFRX1 \CACHE_reg[6][11]  ( .D(n2722), .CK(clk), .RN(n526), .Q(
        \CACHE[6][11] ), .QN(n1482) );
  DFFRX1 \CACHE_reg[6][10]  ( .D(n2721), .CK(clk), .RN(n529), .Q(
        \CACHE[6][10] ), .QN(n1481) );
  DFFRX1 \CACHE_reg[6][9]  ( .D(n2720), .CK(clk), .RN(n532), .Q(\CACHE[6][9] ), 
        .QN(n1480) );
  DFFRX1 \CACHE_reg[6][8]  ( .D(n2719), .CK(clk), .RN(n534), .Q(\CACHE[6][8] ), 
        .QN(n1479) );
  DFFRX1 \CACHE_reg[6][7]  ( .D(n2718), .CK(clk), .RN(n537), .Q(\CACHE[6][7] ), 
        .QN(n1478) );
  DFFRX1 \CACHE_reg[6][6]  ( .D(n2717), .CK(clk), .RN(n540), .Q(\CACHE[6][6] ), 
        .QN(n1477) );
  DFFRX1 \CACHE_reg[6][5]  ( .D(n2716), .CK(clk), .RN(n3022), .Q(\CACHE[6][5] ), .QN(n1476) );
  DFFRX1 \CACHE_reg[6][4]  ( .D(n2715), .CK(clk), .RN(n3058), .Q(\CACHE[6][4] ), .QN(n1475) );
  DFFRX1 \CACHE_reg[6][3]  ( .D(n2714), .CK(clk), .RN(n3025), .Q(\CACHE[6][3] ), .QN(n1474) );
  DFFRX1 \CACHE_reg[6][2]  ( .D(n2713), .CK(clk), .RN(n3028), .Q(\CACHE[6][2] ), .QN(n1473) );
  DFFRX1 \CACHE_reg[6][1]  ( .D(n2712), .CK(clk), .RN(n3039), .Q(\CACHE[6][1] ), .QN(n1472) );
  DFFRX1 \CACHE_reg[6][0]  ( .D(n2711), .CK(clk), .RN(n3030), .Q(\CACHE[6][0] ), .QN(n1471) );
  DFFRX1 \CACHE_reg[2][154]  ( .D(n2245), .CK(clk), .RN(n3057), .Q(
        \CACHE[2][154] ), .QN(n1005) );
  DFFRX1 \CACHE_reg[2][153]  ( .D(n2244), .CK(clk), .RN(n3057), .Q(
        \CACHE[2][153] ), .QN(n1004) );
  DFFRX1 \CACHE_reg[2][152]  ( .D(n2243), .CK(clk), .RN(n3056), .Q(
        \CACHE[2][152] ), .QN(n1003) );
  DFFRX1 \CACHE_reg[2][151]  ( .D(n2242), .CK(clk), .RN(n3040), .Q(
        \CACHE[2][151] ), .QN(n1002) );
  DFFRX1 \CACHE_reg[2][150]  ( .D(n2241), .CK(clk), .RN(n3041), .Q(
        \CACHE[2][150] ), .QN(n1001) );
  DFFRX1 \CACHE_reg[2][149]  ( .D(n2240), .CK(clk), .RN(n3041), .Q(
        \CACHE[2][149] ), .QN(n1000) );
  DFFRX1 \CACHE_reg[2][148]  ( .D(n2239), .CK(clk), .RN(n3042), .Q(
        \CACHE[2][148] ), .QN(n999) );
  DFFRX1 \CACHE_reg[2][147]  ( .D(n2238), .CK(clk), .RN(n3043), .Q(
        \CACHE[2][147] ), .QN(n998) );
  DFFRX1 \CACHE_reg[2][146]  ( .D(n2237), .CK(clk), .RN(n3043), .Q(
        \CACHE[2][146] ), .QN(n997) );
  DFFRX1 \CACHE_reg[2][145]  ( .D(n2236), .CK(clk), .RN(n3044), .Q(
        \CACHE[2][145] ), .QN(n996) );
  DFFRX1 \CACHE_reg[2][144]  ( .D(n2235), .CK(clk), .RN(n3045), .Q(
        \CACHE[2][144] ), .QN(n995) );
  DFFRX1 \CACHE_reg[2][143]  ( .D(n2234), .CK(clk), .RN(n3045), .Q(
        \CACHE[2][143] ), .QN(n994) );
  DFFRX1 \CACHE_reg[2][142]  ( .D(n2233), .CK(clk), .RN(n3046), .Q(
        \CACHE[2][142] ), .QN(n993) );
  DFFRX1 \CACHE_reg[2][141]  ( .D(n2232), .CK(clk), .RN(n3047), .Q(
        \CACHE[2][141] ), .QN(n992) );
  DFFRX1 \CACHE_reg[2][140]  ( .D(n2231), .CK(clk), .RN(n3047), .Q(
        \CACHE[2][140] ), .QN(n991) );
  DFFRX1 \CACHE_reg[2][139]  ( .D(n2230), .CK(clk), .RN(n3048), .Q(
        \CACHE[2][139] ), .QN(n990) );
  DFFRX1 \CACHE_reg[2][138]  ( .D(n2229), .CK(clk), .RN(n3049), .Q(
        \CACHE[2][138] ), .QN(n989) );
  DFFRX1 \CACHE_reg[2][137]  ( .D(n2228), .CK(clk), .RN(n3049), .Q(
        \CACHE[2][137] ), .QN(n988) );
  DFFRX1 \CACHE_reg[2][136]  ( .D(n2227), .CK(clk), .RN(n3050), .Q(
        \CACHE[2][136] ), .QN(n987) );
  DFFRX1 \CACHE_reg[2][135]  ( .D(n2226), .CK(clk), .RN(n3051), .Q(
        \CACHE[2][135] ), .QN(n986) );
  DFFRX1 \CACHE_reg[2][134]  ( .D(n2225), .CK(clk), .RN(n3051), .Q(
        \CACHE[2][134] ), .QN(n985) );
  DFFRX1 \CACHE_reg[2][133]  ( .D(n2224), .CK(clk), .RN(n3052), .Q(
        \CACHE[2][133] ), .QN(n984) );
  DFFRX1 \CACHE_reg[2][132]  ( .D(n2223), .CK(clk), .RN(n3053), .Q(
        \CACHE[2][132] ), .QN(n983) );
  DFFRX1 \CACHE_reg[2][131]  ( .D(n2222), .CK(clk), .RN(n3053), .Q(
        \CACHE[2][131] ), .QN(n982) );
  DFFRX1 \CACHE_reg[2][130]  ( .D(n2221), .CK(clk), .RN(n3054), .Q(
        \CACHE[2][130] ), .QN(n981) );
  DFFRX1 \CACHE_reg[2][129]  ( .D(n2220), .CK(clk), .RN(n3055), .Q(
        \CACHE[2][129] ), .QN(n980) );
  DFFRX1 \CACHE_reg[2][128]  ( .D(n2219), .CK(clk), .RN(n3055), .Q(
        \CACHE[2][128] ), .QN(n979) );
  DFFRX1 \CACHE_reg[2][127]  ( .D(n2218), .CK(clk), .RN(n478), .Q(
        \CACHE[2][127] ), .QN(n978) );
  DFFRX1 \CACHE_reg[2][126]  ( .D(n2217), .CK(clk), .RN(n481), .Q(
        \CACHE[2][126] ), .QN(n977) );
  DFFRX1 \CACHE_reg[2][125]  ( .D(n2216), .CK(clk), .RN(n483), .Q(
        \CACHE[2][125] ), .QN(n976) );
  DFFRX1 \CACHE_reg[2][124]  ( .D(n2215), .CK(clk), .RN(n486), .Q(
        \CACHE[2][124] ), .QN(n975) );
  DFFRX1 \CACHE_reg[2][123]  ( .D(n2214), .CK(clk), .RN(n489), .Q(
        \CACHE[2][123] ), .QN(n974) );
  DFFRX1 \CACHE_reg[2][122]  ( .D(n2213), .CK(clk), .RN(n491), .Q(
        \CACHE[2][122] ), .QN(n973) );
  DFFRX1 \CACHE_reg[2][121]  ( .D(n2212), .CK(clk), .RN(n494), .Q(
        \CACHE[2][121] ), .QN(n972) );
  DFFRX1 \CACHE_reg[2][120]  ( .D(n2211), .CK(clk), .RN(n497), .Q(
        \CACHE[2][120] ), .QN(n971) );
  DFFRX1 \CACHE_reg[2][119]  ( .D(n2210), .CK(clk), .RN(n499), .Q(
        \CACHE[2][119] ), .QN(n970) );
  DFFRX1 \CACHE_reg[2][118]  ( .D(n2209), .CK(clk), .RN(n502), .Q(
        \CACHE[2][118] ), .QN(n969) );
  DFFRX1 \CACHE_reg[2][117]  ( .D(n2208), .CK(clk), .RN(n505), .Q(
        \CACHE[2][117] ), .QN(n968) );
  DFFRX1 \CACHE_reg[2][116]  ( .D(n2207), .CK(clk), .RN(n507), .Q(
        \CACHE[2][116] ), .QN(n967) );
  DFFRX1 \CACHE_reg[2][115]  ( .D(n2206), .CK(clk), .RN(n510), .Q(
        \CACHE[2][115] ), .QN(n966) );
  DFFRX1 \CACHE_reg[2][114]  ( .D(n2205), .CK(clk), .RN(n3033), .Q(
        \CACHE[2][114] ), .QN(n965) );
  DFFRX1 \CACHE_reg[2][113]  ( .D(n2204), .CK(clk), .RN(n513), .Q(
        \CACHE[2][113] ), .QN(n964) );
  DFFRX1 \CACHE_reg[2][112]  ( .D(n2203), .CK(clk), .RN(n515), .Q(
        \CACHE[2][112] ), .QN(n963) );
  DFFRX1 \CACHE_reg[2][111]  ( .D(n2202), .CK(clk), .RN(n518), .Q(
        \CACHE[2][111] ), .QN(n962) );
  DFFRX1 \CACHE_reg[2][110]  ( .D(n2201), .CK(clk), .RN(n521), .Q(
        \CACHE[2][110] ), .QN(n961) );
  DFFRX1 \CACHE_reg[2][109]  ( .D(n2200), .CK(clk), .RN(n523), .Q(
        \CACHE[2][109] ), .QN(n960) );
  DFFRX1 \CACHE_reg[2][108]  ( .D(n2199), .CK(clk), .RN(n526), .Q(
        \CACHE[2][108] ), .QN(n959) );
  DFFRX1 \CACHE_reg[2][107]  ( .D(n2198), .CK(clk), .RN(n529), .Q(
        \CACHE[2][107] ), .QN(n958) );
  DFFRX1 \CACHE_reg[2][106]  ( .D(n2197), .CK(clk), .RN(n531), .Q(
        \CACHE[2][106] ), .QN(n957) );
  DFFRX1 \CACHE_reg[2][105]  ( .D(n2196), .CK(clk), .RN(n534), .Q(
        \CACHE[2][105] ), .QN(n956) );
  DFFRX1 \CACHE_reg[2][104]  ( .D(n2195), .CK(clk), .RN(n537), .Q(
        \CACHE[2][104] ), .QN(n955) );
  DFFRX1 \CACHE_reg[2][103]  ( .D(n2194), .CK(clk), .RN(n539), .Q(
        \CACHE[2][103] ), .QN(n954) );
  DFFRX1 \CACHE_reg[2][102]  ( .D(n2193), .CK(clk), .RN(n3022), .Q(
        \CACHE[2][102] ), .QN(n953) );
  DFFRX1 \CACHE_reg[2][101]  ( .D(n2192), .CK(clk), .RN(n3025), .Q(
        \CACHE[2][101] ), .QN(n952) );
  DFFRX1 \CACHE_reg[2][100]  ( .D(n2191), .CK(clk), .RN(n3034), .Q(
        \CACHE[2][100] ), .QN(n951) );
  DFFRX1 \CACHE_reg[2][99]  ( .D(n2190), .CK(clk), .RN(n3027), .Q(
        \CACHE[2][99] ), .QN(n950) );
  DFFRX1 \CACHE_reg[2][98]  ( .D(n2189), .CK(clk), .RN(n3030), .Q(
        \CACHE[2][98] ), .QN(n949) );
  DFFRX1 \CACHE_reg[2][97]  ( .D(n2188), .CK(clk), .RN(n3035), .Q(
        \CACHE[2][97] ), .QN(n948) );
  DFFRX1 \CACHE_reg[2][96]  ( .D(n2187), .CK(clk), .RN(n3033), .Q(
        \CACHE[2][96] ), .QN(n947) );
  DFFRX1 \CACHE_reg[2][95]  ( .D(n2186), .CK(clk), .RN(n477), .Q(
        \CACHE[2][95] ), .QN(n946) );
  DFFRX1 \CACHE_reg[2][94]  ( .D(n2185), .CK(clk), .RN(n480), .Q(
        \CACHE[2][94] ), .QN(n945) );
  DFFRX1 \CACHE_reg[2][93]  ( .D(n2184), .CK(clk), .RN(n483), .Q(
        \CACHE[2][93] ), .QN(n944) );
  DFFRX1 \CACHE_reg[2][92]  ( .D(n2183), .CK(clk), .RN(n485), .Q(
        \CACHE[2][92] ), .QN(n943) );
  DFFRX1 \CACHE_reg[2][91]  ( .D(n2182), .CK(clk), .RN(n488), .Q(
        \CACHE[2][91] ), .QN(n942) );
  DFFRX1 \CACHE_reg[2][90]  ( .D(n2181), .CK(clk), .RN(n491), .Q(
        \CACHE[2][90] ), .QN(n941) );
  DFFRX1 \CACHE_reg[2][89]  ( .D(n2180), .CK(clk), .RN(n493), .Q(
        \CACHE[2][89] ), .QN(n940) );
  DFFRX1 \CACHE_reg[2][88]  ( .D(n2179), .CK(clk), .RN(n496), .Q(
        \CACHE[2][88] ), .QN(n939) );
  DFFRX1 \CACHE_reg[2][87]  ( .D(n2178), .CK(clk), .RN(n499), .Q(
        \CACHE[2][87] ), .QN(n938) );
  DFFRX1 \CACHE_reg[2][86]  ( .D(n2177), .CK(clk), .RN(n501), .Q(
        \CACHE[2][86] ), .QN(n937) );
  DFFRX1 \CACHE_reg[2][85]  ( .D(n2176), .CK(clk), .RN(n504), .Q(
        \CACHE[2][85] ), .QN(n936) );
  DFFRX1 \CACHE_reg[2][84]  ( .D(n2175), .CK(clk), .RN(n507), .Q(
        \CACHE[2][84] ), .QN(n935) );
  DFFRX1 \CACHE_reg[2][83]  ( .D(n2174), .CK(clk), .RN(n509), .Q(
        \CACHE[2][83] ), .QN(n934) );
  DFFRX1 \CACHE_reg[2][82]  ( .D(n2173), .CK(clk), .RN(n3035), .Q(
        \CACHE[2][82] ), .QN(n933) );
  DFFRX1 \CACHE_reg[2][81]  ( .D(n2172), .CK(clk), .RN(n512), .Q(
        \CACHE[2][81] ), .QN(n932) );
  DFFRX1 \CACHE_reg[2][80]  ( .D(n2171), .CK(clk), .RN(n515), .Q(
        \CACHE[2][80] ), .QN(n931) );
  DFFRX1 \CACHE_reg[2][79]  ( .D(n2170), .CK(clk), .RN(n517), .Q(
        \CACHE[2][79] ), .QN(n930) );
  DFFRX1 \CACHE_reg[2][78]  ( .D(n2169), .CK(clk), .RN(n520), .Q(
        \CACHE[2][78] ), .QN(n929) );
  DFFRX1 \CACHE_reg[2][77]  ( .D(n2168), .CK(clk), .RN(n523), .Q(
        \CACHE[2][77] ), .QN(n928) );
  DFFRX1 \CACHE_reg[2][76]  ( .D(n2167), .CK(clk), .RN(n525), .Q(
        \CACHE[2][76] ), .QN(n927) );
  DFFRX1 \CACHE_reg[2][75]  ( .D(n2166), .CK(clk), .RN(n528), .Q(
        \CACHE[2][75] ), .QN(n926) );
  DFFRX1 \CACHE_reg[2][74]  ( .D(n2165), .CK(clk), .RN(n531), .Q(
        \CACHE[2][74] ), .QN(n925) );
  DFFRX1 \CACHE_reg[2][73]  ( .D(n2164), .CK(clk), .RN(n533), .Q(
        \CACHE[2][73] ), .QN(n924) );
  DFFRX1 \CACHE_reg[2][72]  ( .D(n2163), .CK(clk), .RN(n536), .Q(
        \CACHE[2][72] ), .QN(n923) );
  DFFRX1 \CACHE_reg[2][71]  ( .D(n2162), .CK(clk), .RN(n539), .Q(
        \CACHE[2][71] ), .QN(n922) );
  DFFRX1 \CACHE_reg[2][70]  ( .D(n2161), .CK(clk), .RN(n3020), .Q(
        \CACHE[2][70] ), .QN(n921) );
  DFFRX1 \CACHE_reg[2][69]  ( .D(n2160), .CK(clk), .RN(n3024), .Q(
        \CACHE[2][69] ), .QN(n920) );
  DFFRX1 \CACHE_reg[2][68]  ( .D(n2159), .CK(clk), .RN(n3036), .Q(
        \CACHE[2][68] ), .QN(n919) );
  DFFRX1 \CACHE_reg[2][67]  ( .D(n2158), .CK(clk), .RN(n3027), .Q(
        \CACHE[2][67] ), .QN(n918) );
  DFFRX1 \CACHE_reg[2][66]  ( .D(n2157), .CK(clk), .RN(n3029), .Q(
        \CACHE[2][66] ), .QN(n917) );
  DFFRX1 \CACHE_reg[2][65]  ( .D(n2156), .CK(clk), .RN(n3037), .Q(
        \CACHE[2][65] ), .QN(n916) );
  DFFRX1 \CACHE_reg[2][64]  ( .D(n2155), .CK(clk), .RN(n3032), .Q(
        \CACHE[2][64] ), .QN(n915) );
  DFFRX1 \CACHE_reg[2][63]  ( .D(n2154), .CK(clk), .RN(n477), .Q(
        \CACHE[2][63] ), .QN(n914) );
  DFFRX1 \CACHE_reg[2][62]  ( .D(n2153), .CK(clk), .RN(n479), .Q(
        \CACHE[2][62] ), .QN(n913) );
  DFFRX1 \CACHE_reg[2][61]  ( .D(n2152), .CK(clk), .RN(n482), .Q(
        \CACHE[2][61] ), .QN(n912) );
  DFFRX1 \CACHE_reg[2][60]  ( .D(n2151), .CK(clk), .RN(n485), .Q(
        \CACHE[2][60] ), .QN(n911) );
  DFFRX1 \CACHE_reg[2][59]  ( .D(n2150), .CK(clk), .RN(n487), .Q(
        \CACHE[2][59] ), .QN(n910) );
  DFFRX1 \CACHE_reg[2][58]  ( .D(n2149), .CK(clk), .RN(n490), .Q(
        \CACHE[2][58] ), .QN(n909) );
  DFFRX1 \CACHE_reg[2][57]  ( .D(n2148), .CK(clk), .RN(n493), .Q(
        \CACHE[2][57] ), .QN(n908) );
  DFFRX1 \CACHE_reg[2][56]  ( .D(n2147), .CK(clk), .RN(n495), .Q(
        \CACHE[2][56] ), .QN(n907) );
  DFFRX1 \CACHE_reg[2][55]  ( .D(n2146), .CK(clk), .RN(n498), .Q(
        \CACHE[2][55] ), .QN(n906) );
  DFFRX1 \CACHE_reg[2][54]  ( .D(n2145), .CK(clk), .RN(n501), .Q(
        \CACHE[2][54] ), .QN(n905) );
  DFFRX1 \CACHE_reg[2][53]  ( .D(n2144), .CK(clk), .RN(n503), .Q(
        \CACHE[2][53] ), .QN(n904) );
  DFFRX1 \CACHE_reg[2][52]  ( .D(n2143), .CK(clk), .RN(n506), .Q(
        \CACHE[2][52] ), .QN(n903) );
  DFFRX1 \CACHE_reg[2][51]  ( .D(n2142), .CK(clk), .RN(n509), .Q(
        \CACHE[2][51] ), .QN(n902) );
  DFFRX1 \CACHE_reg[2][50]  ( .D(n2141), .CK(clk), .RN(n3037), .Q(
        \CACHE[2][50] ), .QN(n901) );
  DFFRX1 \CACHE_reg[2][49]  ( .D(n2140), .CK(clk), .RN(n511), .Q(
        \CACHE[2][49] ), .QN(n900) );
  DFFRX1 \CACHE_reg[2][48]  ( .D(n2139), .CK(clk), .RN(n514), .Q(
        \CACHE[2][48] ), .QN(n899) );
  DFFRX1 \CACHE_reg[2][47]  ( .D(n2138), .CK(clk), .RN(n517), .Q(
        \CACHE[2][47] ), .QN(n898) );
  DFFRX1 \CACHE_reg[2][46]  ( .D(n2137), .CK(clk), .RN(n519), .Q(
        \CACHE[2][46] ), .QN(n897) );
  DFFRX1 \CACHE_reg[2][45]  ( .D(n2136), .CK(clk), .RN(n522), .Q(
        \CACHE[2][45] ), .QN(n896) );
  DFFRX1 \CACHE_reg[2][44]  ( .D(n2135), .CK(clk), .RN(n525), .Q(
        \CACHE[2][44] ), .QN(n895) );
  DFFRX1 \CACHE_reg[2][43]  ( .D(n2134), .CK(clk), .RN(n527), .Q(
        \CACHE[2][43] ), .QN(n894) );
  DFFRX1 \CACHE_reg[2][42]  ( .D(n2133), .CK(clk), .RN(n530), .Q(
        \CACHE[2][42] ), .QN(n893) );
  DFFRX1 \CACHE_reg[2][41]  ( .D(n2132), .CK(clk), .RN(n533), .Q(
        \CACHE[2][41] ), .QN(n892) );
  DFFRX1 \CACHE_reg[2][40]  ( .D(n2131), .CK(clk), .RN(n535), .Q(
        \CACHE[2][40] ), .QN(n891) );
  DFFRX1 \CACHE_reg[2][39]  ( .D(n2130), .CK(clk), .RN(n538), .Q(
        \CACHE[2][39] ), .QN(n890) );
  DFFRX1 \CACHE_reg[2][38]  ( .D(n2129), .CK(clk), .RN(n3020), .Q(
        \CACHE[2][38] ), .QN(n889) );
  DFFRX1 \CACHE_reg[2][37]  ( .D(n2128), .CK(clk), .RN(n3023), .Q(
        \CACHE[2][37] ), .QN(n888) );
  DFFRX1 \CACHE_reg[2][36]  ( .D(n2127), .CK(clk), .RN(n3038), .Q(
        \CACHE[2][36] ), .QN(n887) );
  DFFRX1 \CACHE_reg[2][35]  ( .D(n2126), .CK(clk), .RN(n3026), .Q(
        \CACHE[2][35] ), .QN(n886) );
  DFFRX1 \CACHE_reg[2][34]  ( .D(n2125), .CK(clk), .RN(n3029), .Q(
        \CACHE[2][34] ), .QN(n885) );
  DFFRX1 \CACHE_reg[2][33]  ( .D(n2124), .CK(clk), .RN(n3039), .Q(
        \CACHE[2][33] ), .QN(n884) );
  DFFRX1 \CACHE_reg[2][32]  ( .D(n2123), .CK(clk), .RN(n3031), .Q(
        \CACHE[2][32] ), .QN(n883) );
  DFFRX1 \CACHE_reg[2][31]  ( .D(n2122), .CK(clk), .RN(n476), .Q(
        \CACHE[2][31] ), .QN(n882) );
  DFFRX1 \CACHE_reg[2][30]  ( .D(n2121), .CK(clk), .RN(n479), .Q(
        \CACHE[2][30] ), .QN(n881) );
  DFFRX1 \CACHE_reg[2][29]  ( .D(n2120), .CK(clk), .RN(n481), .Q(
        \CACHE[2][29] ), .QN(n880) );
  DFFRX1 \CACHE_reg[2][28]  ( .D(n2119), .CK(clk), .RN(n484), .Q(
        \CACHE[2][28] ), .QN(n879) );
  DFFRX1 \CACHE_reg[2][27]  ( .D(n2118), .CK(clk), .RN(n487), .Q(
        \CACHE[2][27] ), .QN(n878) );
  DFFRX1 \CACHE_reg[2][26]  ( .D(n2117), .CK(clk), .RN(n489), .Q(
        \CACHE[2][26] ), .QN(n877) );
  DFFRX1 \CACHE_reg[2][25]  ( .D(n2116), .CK(clk), .RN(n492), .Q(
        \CACHE[2][25] ), .QN(n876) );
  DFFRX1 \CACHE_reg[2][24]  ( .D(n2115), .CK(clk), .RN(n495), .Q(
        \CACHE[2][24] ), .QN(n875) );
  DFFRX1 \CACHE_reg[2][23]  ( .D(n2114), .CK(clk), .RN(n497), .Q(
        \CACHE[2][23] ), .QN(n874) );
  DFFRX1 \CACHE_reg[2][22]  ( .D(n2113), .CK(clk), .RN(n500), .Q(
        \CACHE[2][22] ), .QN(n873) );
  DFFRX1 \CACHE_reg[2][21]  ( .D(n2112), .CK(clk), .RN(n503), .Q(
        \CACHE[2][21] ), .QN(n872) );
  DFFRX1 \CACHE_reg[2][20]  ( .D(n2111), .CK(clk), .RN(n505), .Q(
        \CACHE[2][20] ), .QN(n871) );
  DFFRX1 \CACHE_reg[2][19]  ( .D(n2110), .CK(clk), .RN(n508), .Q(
        \CACHE[2][19] ), .QN(n870) );
  DFFRX1 \CACHE_reg[2][18]  ( .D(n2109), .CK(clk), .RN(n3059), .Q(
        \CACHE[2][18] ), .QN(n869) );
  DFFRX1 \CACHE_reg[2][17]  ( .D(n2108), .CK(clk), .RN(n511), .Q(
        \CACHE[2][17] ), .QN(n868) );
  DFFRX1 \CACHE_reg[2][16]  ( .D(n2107), .CK(clk), .RN(n513), .Q(
        \CACHE[2][16] ), .QN(n867) );
  DFFRX1 \CACHE_reg[2][15]  ( .D(n2106), .CK(clk), .RN(n516), .Q(
        \CACHE[2][15] ), .QN(n866) );
  DFFRX1 \CACHE_reg[2][14]  ( .D(n2105), .CK(clk), .RN(n519), .Q(
        \CACHE[2][14] ), .QN(n865) );
  DFFRX1 \CACHE_reg[2][13]  ( .D(n2104), .CK(clk), .RN(n521), .Q(
        \CACHE[2][13] ), .QN(n864) );
  DFFRX1 \CACHE_reg[2][12]  ( .D(n2103), .CK(clk), .RN(n524), .Q(
        \CACHE[2][12] ), .QN(n863) );
  DFFRX1 \CACHE_reg[2][11]  ( .D(n2102), .CK(clk), .RN(n527), .Q(
        \CACHE[2][11] ), .QN(n862) );
  DFFRX1 \CACHE_reg[2][10]  ( .D(n2101), .CK(clk), .RN(n529), .Q(
        \CACHE[2][10] ), .QN(n861) );
  DFFRX1 \CACHE_reg[2][9]  ( .D(n2100), .CK(clk), .RN(n532), .Q(\CACHE[2][9] ), 
        .QN(n860) );
  DFFRX1 \CACHE_reg[2][8]  ( .D(n2099), .CK(clk), .RN(n535), .Q(\CACHE[2][8] ), 
        .QN(n859) );
  DFFRX1 \CACHE_reg[2][7]  ( .D(n2098), .CK(clk), .RN(n537), .Q(\CACHE[2][7] ), 
        .QN(n858) );
  DFFRX1 \CACHE_reg[2][6]  ( .D(n2097), .CK(clk), .RN(n540), .Q(\CACHE[2][6] ), 
        .QN(n857) );
  DFFRX1 \CACHE_reg[2][5]  ( .D(n2096), .CK(clk), .RN(n3023), .Q(\CACHE[2][5] ), .QN(n856) );
  DFFRX1 \CACHE_reg[2][4]  ( .D(n2095), .CK(clk), .RN(n3058), .Q(\CACHE[2][4] ), .QN(n855) );
  DFFRX1 \CACHE_reg[2][3]  ( .D(n2094), .CK(clk), .RN(n3025), .Q(\CACHE[2][3] ), .QN(n854) );
  DFFRX1 \CACHE_reg[2][2]  ( .D(n2093), .CK(clk), .RN(n3028), .Q(\CACHE[2][2] ), .QN(n853) );
  DFFRX1 \CACHE_reg[2][1]  ( .D(n2092), .CK(clk), .RN(n3039), .Q(\CACHE[2][1] ), .QN(n852) );
  DFFRX1 \CACHE_reg[2][0]  ( .D(n2091), .CK(clk), .RN(n3031), .Q(\CACHE[2][0] ), .QN(n851) );
  NOR3X6 U3 ( .A(proc_addr[0]), .B(proc_addr[1]), .C(n3742), .Y(n3760) );
  NOR3X6 U4 ( .A(n3575), .B(proc_addr[1]), .C(n3742), .Y(n3757) );
  NOR3X6 U5 ( .A(n3576), .B(proc_addr[0]), .C(n3742), .Y(n3753) );
  AND2X2 U6 ( .A(n3767), .B(mem_ready), .Y(n3744) );
  OR2X1 U7 ( .A(n3768), .B(n475), .Y(n1) );
  AOI22X1 U8 ( .A0(N59), .A1(n415), .B0(proc_addr[5]), .B1(mem_read), .Y(n2)
         );
  AOI22X1 U9 ( .A0(N58), .A1(n415), .B0(proc_addr[6]), .B1(mem_read), .Y(n3)
         );
  AOI22X1 U10 ( .A0(N57), .A1(n415), .B0(proc_addr[7]), .B1(mem_read), .Y(n4)
         );
  AOI22X1 U11 ( .A0(N56), .A1(n416), .B0(proc_addr[8]), .B1(mem_read), .Y(n5)
         );
  AOI22X1 U12 ( .A0(N55), .A1(n417), .B0(proc_addr[9]), .B1(mem_read), .Y(n6)
         );
  AOI22X1 U13 ( .A0(N54), .A1(mem_write), .B0(proc_addr[10]), .B1(mem_read), 
        .Y(n7) );
  AOI22X1 U14 ( .A0(N53), .A1(n413), .B0(proc_addr[11]), .B1(mem_read), .Y(n8)
         );
  AOI22X1 U15 ( .A0(N52), .A1(n413), .B0(proc_addr[12]), .B1(mem_read), .Y(n9)
         );
  AOI22X1 U16 ( .A0(N51), .A1(n416), .B0(proc_addr[13]), .B1(mem_read), .Y(n10) );
  AOI22X1 U17 ( .A0(N50), .A1(mem_write), .B0(proc_addr[14]), .B1(mem_read), 
        .Y(n11) );
  AOI22X1 U18 ( .A0(N49), .A1(n413), .B0(proc_addr[15]), .B1(mem_read), .Y(n12) );
  AOI22X1 U19 ( .A0(N48), .A1(n416), .B0(proc_addr[16]), .B1(mem_read), .Y(n13) );
  AOI22X1 U20 ( .A0(N47), .A1(n417), .B0(proc_addr[17]), .B1(mem_read), .Y(n14) );
  AOI22X1 U21 ( .A0(N46), .A1(n319), .B0(proc_addr[18]), .B1(mem_read), .Y(n15) );
  AOI22X1 U22 ( .A0(N45), .A1(mem_write), .B0(proc_addr[19]), .B1(mem_read), 
        .Y(n16) );
  AOI22X1 U23 ( .A0(N44), .A1(n417), .B0(proc_addr[20]), .B1(mem_read), .Y(n17) );
  AOI22X1 U24 ( .A0(N43), .A1(n413), .B0(proc_addr[21]), .B1(mem_read), .Y(n18) );
  AOI22X1 U25 ( .A0(N42), .A1(mem_write), .B0(proc_addr[22]), .B1(mem_read), 
        .Y(n19) );
  AOI22X1 U26 ( .A0(N41), .A1(mem_write), .B0(proc_addr[23]), .B1(mem_read), 
        .Y(n20) );
  AOI22X1 U27 ( .A0(N40), .A1(mem_write), .B0(proc_addr[24]), .B1(mem_read), 
        .Y(n21) );
  AOI22X1 U28 ( .A0(N39), .A1(n415), .B0(proc_addr[25]), .B1(mem_read), .Y(n22) );
  AOI22X1 U29 ( .A0(N38), .A1(n415), .B0(proc_addr[26]), .B1(mem_read), .Y(n23) );
  AOI22X1 U30 ( .A0(N37), .A1(n415), .B0(proc_addr[27]), .B1(mem_read), .Y(n24) );
  AOI22X1 U31 ( .A0(N36), .A1(n415), .B0(proc_addr[28]), .B1(mem_read), .Y(n25) );
  AOI22X1 U32 ( .A0(N35), .A1(n415), .B0(proc_addr[29]), .B1(mem_read), .Y(n26) );
  OR2X1 U33 ( .A(n3572), .B(n402), .Y(n27) );
  OR2X1 U34 ( .A(n3517), .B(n405), .Y(n28) );
  OR2X1 U35 ( .A(n3462), .B(n406), .Y(n29) );
  OR2X1 U36 ( .A(n3447), .B(n407), .Y(n30) );
  OR2X1 U37 ( .A(n3442), .B(n408), .Y(n31) );
  OR2X1 U38 ( .A(n3437), .B(n408), .Y(n32) );
  OR2X1 U39 ( .A(n3432), .B(n409), .Y(n33) );
  OR2X1 U40 ( .A(n3427), .B(n410), .Y(n34) );
  OR2X1 U41 ( .A(n3422), .B(n411), .Y(n35) );
  OR2X1 U42 ( .A(n3416), .B(n412), .Y(n36) );
  OR2X1 U43 ( .A(n3567), .B(n402), .Y(n37) );
  OR2X1 U44 ( .A(n3562), .B(n403), .Y(n38) );
  OR2X1 U45 ( .A(n3557), .B(n404), .Y(n39) );
  OR2X1 U46 ( .A(n3552), .B(n404), .Y(n40) );
  OR2X1 U47 ( .A(n3547), .B(n404), .Y(n41) );
  OR2X1 U48 ( .A(n3542), .B(n404), .Y(n42) );
  OR2X1 U49 ( .A(n3537), .B(n404), .Y(n43) );
  OR2X1 U50 ( .A(n3532), .B(n405), .Y(n44) );
  OR2X1 U51 ( .A(n3527), .B(n405), .Y(n45) );
  OR2X1 U52 ( .A(n3522), .B(n405), .Y(n46) );
  OR2X1 U53 ( .A(n3512), .B(n405), .Y(n47) );
  OR2X1 U54 ( .A(n3507), .B(n405), .Y(n48) );
  OR2X1 U55 ( .A(n3502), .B(n405), .Y(n49) );
  OR2X1 U56 ( .A(n3497), .B(n405), .Y(n50) );
  OR2X1 U57 ( .A(n3492), .B(n405), .Y(n51) );
  OR2X1 U58 ( .A(n3487), .B(n405), .Y(n52) );
  OR2X1 U59 ( .A(n3482), .B(n405), .Y(n53) );
  OR2X1 U60 ( .A(n3477), .B(n405), .Y(n54) );
  OR2X1 U61 ( .A(n3472), .B(n406), .Y(n55) );
  OR2X1 U62 ( .A(n3467), .B(n406), .Y(n56) );
  OR2X1 U63 ( .A(n3457), .B(n406), .Y(n57) );
  OR2X1 U64 ( .A(n3452), .B(n406), .Y(n58) );
  OR2X1 U65 ( .A(n3570), .B(n406), .Y(n59) );
  OR2X1 U66 ( .A(n3515), .B(n406), .Y(n60) );
  OR2X1 U67 ( .A(n3460), .B(n406), .Y(n61) );
  OR2X1 U68 ( .A(n3445), .B(n406), .Y(n62) );
  OR2X1 U69 ( .A(n3440), .B(n406), .Y(n63) );
  OR2X1 U70 ( .A(n3435), .B(n406), .Y(n64) );
  OR2X1 U71 ( .A(n3430), .B(n406), .Y(n65) );
  OR2X1 U72 ( .A(n3425), .B(n407), .Y(n66) );
  OR2X1 U73 ( .A(n3420), .B(n407), .Y(n67) );
  OR2X1 U74 ( .A(n3414), .B(n407), .Y(n68) );
  OR2X1 U75 ( .A(n3565), .B(n407), .Y(n69) );
  OR2X1 U76 ( .A(n3560), .B(n407), .Y(n70) );
  OR2X1 U77 ( .A(n3555), .B(n407), .Y(n71) );
  OR2X1 U78 ( .A(n3550), .B(n407), .Y(n72) );
  OR2X1 U79 ( .A(n3545), .B(n407), .Y(n73) );
  OR2X1 U80 ( .A(n3540), .B(n407), .Y(n74) );
  OR2X1 U81 ( .A(n3535), .B(n407), .Y(n75) );
  OR2X1 U82 ( .A(n3530), .B(n407), .Y(n76) );
  OR2X1 U83 ( .A(n3525), .B(n408), .Y(n77) );
  OR2X1 U84 ( .A(n3520), .B(n408), .Y(n78) );
  OR2X1 U85 ( .A(n3510), .B(n408), .Y(n79) );
  OR2X1 U86 ( .A(n3505), .B(n408), .Y(n80) );
  OR2X1 U87 ( .A(n3500), .B(n408), .Y(n81) );
  OR2X1 U88 ( .A(n3495), .B(n408), .Y(n82) );
  OR2X1 U89 ( .A(n3490), .B(n408), .Y(n83) );
  OR2X1 U90 ( .A(n3485), .B(n408), .Y(n84) );
  OR2X1 U91 ( .A(n3480), .B(n408), .Y(n85) );
  OR2X1 U92 ( .A(n3475), .B(n408), .Y(n86) );
  OR2X1 U93 ( .A(n3470), .B(n409), .Y(n87) );
  OR2X1 U94 ( .A(n3465), .B(n409), .Y(n88) );
  OR2X1 U95 ( .A(n3455), .B(n409), .Y(n89) );
  OR2X1 U96 ( .A(n3450), .B(n409), .Y(n90) );
  OR2X1 U97 ( .A(n3569), .B(n409), .Y(n91) );
  OR2X1 U98 ( .A(n3514), .B(n409), .Y(n92) );
  OR2X1 U99 ( .A(n3459), .B(n409), .Y(n93) );
  OR2X1 U100 ( .A(n3444), .B(n409), .Y(n94) );
  OR2X1 U101 ( .A(n3439), .B(n409), .Y(n95) );
  OR2X1 U102 ( .A(n3434), .B(n409), .Y(n96) );
  OR2X1 U103 ( .A(n3429), .B(n409), .Y(n97) );
  OR2X1 U104 ( .A(n3424), .B(n410), .Y(n98) );
  OR2X1 U105 ( .A(n3419), .B(n410), .Y(n99) );
  OR2X1 U106 ( .A(n3412), .B(n410), .Y(n100) );
  OR2X1 U107 ( .A(n3564), .B(n410), .Y(n101) );
  OR2X1 U108 ( .A(n3559), .B(n410), .Y(n102) );
  OR2X1 U109 ( .A(n3554), .B(n410), .Y(n103) );
  OR2X1 U110 ( .A(n3549), .B(n410), .Y(n104) );
  OR2X1 U111 ( .A(n3544), .B(n410), .Y(n105) );
  OR2X1 U112 ( .A(n3539), .B(n410), .Y(n106) );
  OR2X1 U113 ( .A(n3534), .B(n410), .Y(n107) );
  OR2X1 U114 ( .A(n3529), .B(n410), .Y(n108) );
  OR2X1 U115 ( .A(n3524), .B(n411), .Y(n109) );
  OR2X1 U116 ( .A(n3519), .B(n411), .Y(n110) );
  OR2X1 U117 ( .A(n3509), .B(n411), .Y(n111) );
  OR2X1 U118 ( .A(n3504), .B(n411), .Y(n112) );
  OR2X1 U119 ( .A(n3499), .B(n411), .Y(n113) );
  OR2X1 U120 ( .A(n3494), .B(n411), .Y(n114) );
  OR2X1 U121 ( .A(n3489), .B(n411), .Y(n115) );
  OR2X1 U122 ( .A(n3484), .B(n411), .Y(n116) );
  OR2X1 U123 ( .A(n3479), .B(n411), .Y(n117) );
  OR2X1 U124 ( .A(n3474), .B(n411), .Y(n118) );
  OR2X1 U125 ( .A(n3469), .B(n411), .Y(n119) );
  OR2X1 U126 ( .A(n3464), .B(n412), .Y(n120) );
  OR2X1 U127 ( .A(n3454), .B(n412), .Y(n121) );
  OR2X1 U128 ( .A(n3449), .B(n412), .Y(n122) );
  OR2X1 U129 ( .A(n3573), .B(n412), .Y(n123) );
  OR2X1 U130 ( .A(n3518), .B(n412), .Y(n124) );
  OR2X1 U131 ( .A(n3463), .B(n412), .Y(n125) );
  OR2X1 U132 ( .A(n3448), .B(n412), .Y(n126) );
  OR2X1 U133 ( .A(n3443), .B(n402), .Y(n127) );
  OR2X1 U134 ( .A(n3438), .B(n402), .Y(n128) );
  OR2X1 U135 ( .A(n3433), .B(n402), .Y(n129) );
  OR2X1 U136 ( .A(n3428), .B(n402), .Y(n130) );
  OR2X1 U137 ( .A(n3423), .B(n402), .Y(n131) );
  OR2X1 U138 ( .A(n3418), .B(n402), .Y(n132) );
  OR2X1 U139 ( .A(n3568), .B(n402), .Y(n133) );
  OR2X1 U140 ( .A(n3563), .B(n402), .Y(n134) );
  OR2X1 U141 ( .A(n3558), .B(n402), .Y(n135) );
  OR2X1 U142 ( .A(n3553), .B(n402), .Y(n136) );
  OR2X1 U143 ( .A(n3548), .B(n403), .Y(n137) );
  OR2X1 U144 ( .A(n3543), .B(n403), .Y(n138) );
  OR2X1 U145 ( .A(n3538), .B(n403), .Y(n139) );
  OR2X1 U146 ( .A(n3533), .B(n403), .Y(n140) );
  OR2X1 U147 ( .A(n3528), .B(n403), .Y(n141) );
  OR2X1 U148 ( .A(n3523), .B(n403), .Y(n142) );
  OR2X1 U149 ( .A(n3513), .B(n403), .Y(n143) );
  OR2X1 U150 ( .A(n3508), .B(n403), .Y(n144) );
  OR2X1 U151 ( .A(n3503), .B(n403), .Y(n145) );
  OR2X1 U152 ( .A(n3498), .B(n403), .Y(n146) );
  OR2X1 U153 ( .A(n3493), .B(n403), .Y(n147) );
  OR2X1 U154 ( .A(n3488), .B(n404), .Y(n148) );
  OR2X1 U155 ( .A(n3483), .B(n404), .Y(n149) );
  OR2X1 U156 ( .A(n3478), .B(n404), .Y(n150) );
  OR2X1 U157 ( .A(n3473), .B(n404), .Y(n151) );
  OR2X1 U158 ( .A(n3468), .B(n404), .Y(n152) );
  OR2X1 U159 ( .A(n3458), .B(n404), .Y(n153) );
  OR2X1 U160 ( .A(n3453), .B(n404), .Y(n154) );
  OR2X1 U161 ( .A(n3768), .B(n437), .Y(n155) );
  OR2X1 U162 ( .A(n3768), .B(n462), .Y(n156) );
  NAND3X6 U163 ( .A(n3575), .B(n3576), .C(n3574), .Y(n157) );
  AND2X2 U164 ( .A(n3574), .B(n3575), .Y(n158) );
  AND2X2 U165 ( .A(n3574), .B(n3576), .Y(n159) );
  AOI22X2 U166 ( .A0(proc_addr[29]), .A1(n394), .B0(n316), .B1(N35), .Y(n3580)
         );
  AOI22X2 U167 ( .A0(proc_addr[28]), .A1(n394), .B0(n316), .B1(N36), .Y(n3581)
         );
  AOI22X2 U168 ( .A0(proc_addr[27]), .A1(n394), .B0(n316), .B1(N37), .Y(n3582)
         );
  AOI22X2 U169 ( .A0(proc_addr[26]), .A1(n394), .B0(n316), .B1(N38), .Y(n3583)
         );
  AOI22X2 U170 ( .A0(proc_addr[25]), .A1(n394), .B0(n316), .B1(N39), .Y(n3584)
         );
  AOI22X2 U171 ( .A0(proc_addr[24]), .A1(n394), .B0(n316), .B1(N40), .Y(n3585)
         );
  AOI22X2 U172 ( .A0(proc_addr[23]), .A1(n394), .B0(n316), .B1(N41), .Y(n3586)
         );
  AOI22X2 U173 ( .A0(proc_addr[22]), .A1(n394), .B0(n316), .B1(N42), .Y(n3587)
         );
  AOI22X2 U174 ( .A0(proc_addr[21]), .A1(n394), .B0(n316), .B1(N43), .Y(n3588)
         );
  AOI22X2 U175 ( .A0(proc_addr[20]), .A1(n394), .B0(n316), .B1(N44), .Y(n3589)
         );
  AOI22X2 U176 ( .A0(proc_addr[19]), .A1(n394), .B0(n316), .B1(N45), .Y(n3590)
         );
  AOI22X2 U177 ( .A0(proc_addr[18]), .A1(n394), .B0(n316), .B1(N46), .Y(n3591)
         );
  AOI22X2 U178 ( .A0(proc_addr[17]), .A1(n401), .B0(n316), .B1(N47), .Y(n3592)
         );
  AOI22X2 U179 ( .A0(proc_addr[16]), .A1(n399), .B0(n316), .B1(N48), .Y(n3593)
         );
  AOI22X2 U180 ( .A0(proc_addr[15]), .A1(n396), .B0(n316), .B1(N49), .Y(n3594)
         );
  AOI22X2 U181 ( .A0(proc_addr[14]), .A1(n398), .B0(n316), .B1(N50), .Y(n3595)
         );
  AOI22X2 U182 ( .A0(proc_addr[13]), .A1(n397), .B0(n316), .B1(N51), .Y(n3596)
         );
  AOI22X2 U183 ( .A0(proc_addr[12]), .A1(n395), .B0(n316), .B1(N52), .Y(n3597)
         );
  AOI22X2 U184 ( .A0(proc_addr[11]), .A1(n400), .B0(n316), .B1(N53), .Y(n3598)
         );
  AOI22X2 U185 ( .A0(proc_addr[7]), .A1(n394), .B0(n316), .B1(N57), .Y(n3602)
         );
  AOI22X2 U186 ( .A0(proc_addr[6]), .A1(n401), .B0(n316), .B1(N58), .Y(n3603)
         );
  AOI22X2 U187 ( .A0(proc_addr[5]), .A1(n400), .B0(n3745), .B1(N59), .Y(n3604)
         );
  AOI222X4 U188 ( .A0(mem_rdata[127]), .A1(n397), .B0(n3748), .B1(N60), .C0(
        proc_wdata[31]), .C1(n3749), .Y(n3605) );
  AOI222X4 U189 ( .A0(mem_rdata[126]), .A1(n395), .B0(n3748), .B1(N61), .C0(
        proc_wdata[30]), .C1(n3749), .Y(n3606) );
  AOI222X4 U190 ( .A0(mem_rdata[125]), .A1(n394), .B0(n3748), .B1(N62), .C0(
        proc_wdata[29]), .C1(n3749), .Y(n3607) );
  AOI222X4 U191 ( .A0(mem_rdata[124]), .A1(n401), .B0(n3748), .B1(N63), .C0(
        proc_wdata[28]), .C1(n3749), .Y(n3608) );
  AOI222X4 U192 ( .A0(mem_rdata[123]), .A1(n399), .B0(n3748), .B1(N64), .C0(
        proc_wdata[27]), .C1(n3749), .Y(n3609) );
  AOI222X4 U193 ( .A0(mem_rdata[122]), .A1(n397), .B0(n3748), .B1(N65), .C0(
        proc_wdata[26]), .C1(n3749), .Y(n3610) );
  AOI222X4 U194 ( .A0(mem_rdata[121]), .A1(n395), .B0(n3748), .B1(N66), .C0(
        proc_wdata[25]), .C1(n3749), .Y(n3611) );
  AOI222X4 U195 ( .A0(mem_rdata[120]), .A1(n3744), .B0(n3748), .B1(N67), .C0(
        proc_wdata[24]), .C1(n3749), .Y(n3612) );
  AOI222X4 U196 ( .A0(mem_rdata[119]), .A1(n3744), .B0(n3748), .B1(N68), .C0(
        proc_wdata[23]), .C1(n3749), .Y(n3613) );
  AOI222X4 U197 ( .A0(mem_rdata[118]), .A1(n3744), .B0(n3748), .B1(N69), .C0(
        proc_wdata[22]), .C1(n3749), .Y(n3614) );
  AOI222X4 U198 ( .A0(mem_rdata[117]), .A1(n3744), .B0(n3748), .B1(N70), .C0(
        proc_wdata[21]), .C1(n3749), .Y(n3615) );
  AOI222X4 U199 ( .A0(mem_rdata[116]), .A1(n395), .B0(n3748), .B1(N71), .C0(
        proc_wdata[20]), .C1(n3749), .Y(n3616) );
  AOI222X4 U200 ( .A0(mem_rdata[115]), .A1(n395), .B0(n3748), .B1(N72), .C0(
        proc_wdata[19]), .C1(n3749), .Y(n3617) );
  AOI222X4 U201 ( .A0(mem_rdata[114]), .A1(n395), .B0(n3748), .B1(N73), .C0(
        proc_wdata[18]), .C1(n3749), .Y(n3618) );
  AOI222X4 U202 ( .A0(mem_rdata[113]), .A1(n395), .B0(n3748), .B1(N74), .C0(
        proc_wdata[17]), .C1(n3749), .Y(n3619) );
  AOI222X4 U203 ( .A0(mem_rdata[112]), .A1(n395), .B0(n3748), .B1(N75), .C0(
        proc_wdata[16]), .C1(n3749), .Y(n3620) );
  AOI222X4 U204 ( .A0(mem_rdata[111]), .A1(n395), .B0(n3748), .B1(N76), .C0(
        proc_wdata[15]), .C1(n3749), .Y(n3621) );
  AOI222X4 U205 ( .A0(mem_rdata[110]), .A1(n395), .B0(n3748), .B1(N77), .C0(
        proc_wdata[14]), .C1(n3749), .Y(n3622) );
  AOI222X4 U206 ( .A0(mem_rdata[109]), .A1(n395), .B0(n3748), .B1(N78), .C0(
        proc_wdata[13]), .C1(n3749), .Y(n3623) );
  AOI222X4 U207 ( .A0(mem_rdata[108]), .A1(n395), .B0(n3748), .B1(N79), .C0(
        proc_wdata[12]), .C1(n3749), .Y(n3624) );
  AOI222X4 U208 ( .A0(mem_rdata[107]), .A1(n395), .B0(n3748), .B1(N80), .C0(
        proc_wdata[11]), .C1(n3749), .Y(n3625) );
  AOI222X4 U209 ( .A0(mem_rdata[106]), .A1(n395), .B0(n3748), .B1(N81), .C0(
        proc_wdata[10]), .C1(n3749), .Y(n3626) );
  AOI222X4 U210 ( .A0(mem_rdata[105]), .A1(n395), .B0(n3748), .B1(N82), .C0(
        proc_wdata[9]), .C1(n3749), .Y(n3627) );
  AOI222X4 U211 ( .A0(mem_rdata[104]), .A1(n395), .B0(n3748), .B1(N83), .C0(
        proc_wdata[8]), .C1(n3749), .Y(n3628) );
  AOI222X4 U212 ( .A0(mem_rdata[103]), .A1(n395), .B0(n3748), .B1(N84), .C0(
        proc_wdata[7]), .C1(n3749), .Y(n3629) );
  AOI222X4 U213 ( .A0(mem_rdata[102]), .A1(n396), .B0(n3748), .B1(N85), .C0(
        proc_wdata[6]), .C1(n3749), .Y(n3630) );
  AOI222X4 U214 ( .A0(mem_rdata[101]), .A1(n396), .B0(n3748), .B1(N86), .C0(
        proc_wdata[5]), .C1(n3749), .Y(n3631) );
  AOI222X4 U215 ( .A0(mem_rdata[100]), .A1(n396), .B0(n3748), .B1(N87), .C0(
        proc_wdata[4]), .C1(n3749), .Y(n3632) );
  AOI222X4 U216 ( .A0(mem_rdata[99]), .A1(n396), .B0(n3748), .B1(N88), .C0(
        proc_wdata[3]), .C1(n3749), .Y(n3633) );
  AOI222X4 U217 ( .A0(mem_rdata[98]), .A1(n396), .B0(n3748), .B1(N89), .C0(
        proc_wdata[2]), .C1(n3749), .Y(n3634) );
  AOI222X4 U218 ( .A0(mem_rdata[97]), .A1(n396), .B0(n3748), .B1(N90), .C0(
        proc_wdata[1]), .C1(n3749), .Y(n3635) );
  AOI222X4 U219 ( .A0(mem_rdata[96]), .A1(n396), .B0(n3748), .B1(N91), .C0(
        proc_wdata[0]), .C1(n3749), .Y(n3636) );
  AOI222X4 U220 ( .A0(n400), .A1(mem_rdata[95]), .B0(proc_wdata[31]), .B1(
        n3753), .C0(N92), .C1(n3754), .Y(n3637) );
  AOI222X4 U221 ( .A0(n398), .A1(mem_rdata[94]), .B0(proc_wdata[30]), .B1(
        n3753), .C0(N93), .C1(n3754), .Y(n3638) );
  AOI222X4 U222 ( .A0(n397), .A1(mem_rdata[93]), .B0(proc_wdata[29]), .B1(
        n3753), .C0(N94), .C1(n3754), .Y(n3639) );
  AOI222X4 U223 ( .A0(n395), .A1(mem_rdata[92]), .B0(proc_wdata[28]), .B1(
        n3753), .C0(N95), .C1(n3754), .Y(n3640) );
  AOI222X4 U224 ( .A0(n400), .A1(mem_rdata[91]), .B0(proc_wdata[27]), .B1(
        n3753), .C0(N96), .C1(n3754), .Y(n3641) );
  AOI222X4 U225 ( .A0(n401), .A1(mem_rdata[90]), .B0(proc_wdata[26]), .B1(
        n3753), .C0(N97), .C1(n3754), .Y(n3642) );
  AOI222X4 U226 ( .A0(n398), .A1(mem_rdata[89]), .B0(proc_wdata[25]), .B1(
        n3753), .C0(N98), .C1(n3754), .Y(n3643) );
  AOI222X4 U227 ( .A0(n3744), .A1(mem_rdata[88]), .B0(proc_wdata[24]), .B1(
        n3753), .C0(N99), .C1(n3754), .Y(n3644) );
  AOI222X4 U228 ( .A0(n401), .A1(mem_rdata[87]), .B0(proc_wdata[23]), .B1(
        n3753), .C0(N100), .C1(n3754), .Y(n3645) );
  AOI222X4 U229 ( .A0(n397), .A1(mem_rdata[86]), .B0(proc_wdata[22]), .B1(
        n3753), .C0(N101), .C1(n3754), .Y(n3646) );
  AOI222X4 U230 ( .A0(n401), .A1(mem_rdata[85]), .B0(proc_wdata[21]), .B1(
        n3753), .C0(N102), .C1(n3754), .Y(n3647) );
  AOI222X4 U231 ( .A0(n401), .A1(mem_rdata[84]), .B0(proc_wdata[20]), .B1(
        n3753), .C0(N103), .C1(n3754), .Y(n3648) );
  AOI222X4 U232 ( .A0(n395), .A1(mem_rdata[83]), .B0(proc_wdata[19]), .B1(
        n3753), .C0(N104), .C1(n3754), .Y(n3649) );
  AOI222X4 U233 ( .A0(n401), .A1(mem_rdata[82]), .B0(proc_wdata[18]), .B1(
        n3753), .C0(N105), .C1(n3754), .Y(n3650) );
  AOI222X4 U234 ( .A0(n401), .A1(mem_rdata[81]), .B0(proc_wdata[17]), .B1(
        n3753), .C0(N106), .C1(n3754), .Y(n3651) );
  AOI222X4 U235 ( .A0(n3744), .A1(mem_rdata[80]), .B0(proc_wdata[16]), .B1(
        n3753), .C0(N107), .C1(n3754), .Y(n3652) );
  AOI222X4 U236 ( .A0(n401), .A1(mem_rdata[79]), .B0(proc_wdata[15]), .B1(
        n3753), .C0(N108), .C1(n3754), .Y(n3653) );
  AOI222X4 U237 ( .A0(n401), .A1(mem_rdata[78]), .B0(proc_wdata[14]), .B1(
        n3753), .C0(N109), .C1(n3754), .Y(n3654) );
  AOI222X4 U238 ( .A0(n396), .A1(mem_rdata[77]), .B0(proc_wdata[13]), .B1(
        n3753), .C0(N110), .C1(n3754), .Y(n3655) );
  AOI222X4 U239 ( .A0(n401), .A1(mem_rdata[76]), .B0(proc_wdata[12]), .B1(
        n3753), .C0(N111), .C1(n3754), .Y(n3656) );
  AOI222X4 U240 ( .A0(n401), .A1(mem_rdata[75]), .B0(proc_wdata[11]), .B1(
        n3753), .C0(N112), .C1(n3754), .Y(n3657) );
  AOI222X4 U241 ( .A0(n400), .A1(mem_rdata[74]), .B0(proc_wdata[10]), .B1(
        n3753), .C0(N113), .C1(n3754), .Y(n3658) );
  AOI222X4 U242 ( .A0(n401), .A1(mem_rdata[73]), .B0(proc_wdata[9]), .B1(n3753), .C0(N114), .C1(n3754), .Y(n3659) );
  AOI222X4 U243 ( .A0(n398), .A1(mem_rdata[72]), .B0(proc_wdata[8]), .B1(n3753), .C0(N115), .C1(n3754), .Y(n3660) );
  AOI222X4 U244 ( .A0(n397), .A1(mem_rdata[71]), .B0(proc_wdata[7]), .B1(n3753), .C0(N116), .C1(n3754), .Y(n3661) );
  AOI222X4 U245 ( .A0(n401), .A1(mem_rdata[70]), .B0(proc_wdata[6]), .B1(n3753), .C0(N117), .C1(n3754), .Y(n3662) );
  AOI222X4 U246 ( .A0(n401), .A1(mem_rdata[69]), .B0(proc_wdata[5]), .B1(n3753), .C0(N118), .C1(n3754), .Y(n3663) );
  AOI222X4 U247 ( .A0(n395), .A1(mem_rdata[68]), .B0(proc_wdata[4]), .B1(n3753), .C0(N119), .C1(n3754), .Y(n3664) );
  AOI222X4 U248 ( .A0(n401), .A1(mem_rdata[67]), .B0(proc_wdata[3]), .B1(n3753), .C0(N120), .C1(n3754), .Y(n3665) );
  AOI222X4 U249 ( .A0(n401), .A1(mem_rdata[66]), .B0(proc_wdata[2]), .B1(n3753), .C0(N121), .C1(n3754), .Y(n3666) );
  AOI222X4 U250 ( .A0(n394), .A1(mem_rdata[65]), .B0(proc_wdata[1]), .B1(n3753), .C0(N122), .C1(n3754), .Y(n3667) );
  AOI222X4 U251 ( .A0(n399), .A1(mem_rdata[64]), .B0(proc_wdata[0]), .B1(n3753), .C0(N123), .C1(n3754), .Y(n3668) );
  AOI222X4 U252 ( .A0(mem_rdata[63]), .A1(n396), .B0(n3756), .B1(N124), .C0(
        n3757), .C1(proc_wdata[31]), .Y(n3669) );
  AOI222X4 U253 ( .A0(mem_rdata[62]), .A1(n396), .B0(n3756), .B1(N125), .C0(
        n3757), .C1(proc_wdata[30]), .Y(n3670) );
  AOI222X4 U254 ( .A0(mem_rdata[61]), .A1(n396), .B0(n3756), .B1(N126), .C0(
        n3757), .C1(proc_wdata[29]), .Y(n3671) );
  AOI222X4 U255 ( .A0(mem_rdata[60]), .A1(n396), .B0(n3756), .B1(N127), .C0(
        n3757), .C1(proc_wdata[28]), .Y(n3672) );
  AOI222X4 U256 ( .A0(mem_rdata[59]), .A1(n396), .B0(n3756), .B1(N128), .C0(
        n3757), .C1(proc_wdata[27]), .Y(n3673) );
  AOI222X4 U257 ( .A0(mem_rdata[58]), .A1(n397), .B0(n3756), .B1(N129), .C0(
        n3757), .C1(proc_wdata[26]), .Y(n3674) );
  AOI222X4 U258 ( .A0(mem_rdata[57]), .A1(n398), .B0(n3756), .B1(N130), .C0(
        n3757), .C1(proc_wdata[25]), .Y(n3675) );
  AOI222X4 U259 ( .A0(mem_rdata[56]), .A1(n396), .B0(n3756), .B1(N131), .C0(
        n3757), .C1(proc_wdata[24]), .Y(n3676) );
  AOI222X4 U260 ( .A0(mem_rdata[55]), .A1(n398), .B0(n3756), .B1(N132), .C0(
        n3757), .C1(proc_wdata[23]), .Y(n3677) );
  AOI222X4 U261 ( .A0(mem_rdata[54]), .A1(n398), .B0(n3756), .B1(N133), .C0(
        n3757), .C1(proc_wdata[22]), .Y(n3678) );
  AOI222X4 U262 ( .A0(mem_rdata[53]), .A1(n397), .B0(n3756), .B1(N134), .C0(
        n3757), .C1(proc_wdata[21]), .Y(n3679) );
  AOI222X4 U263 ( .A0(mem_rdata[52]), .A1(n398), .B0(n3756), .B1(N135), .C0(
        n3757), .C1(proc_wdata[20]), .Y(n3680) );
  AOI222X4 U264 ( .A0(mem_rdata[51]), .A1(n398), .B0(n3756), .B1(N136), .C0(
        n3757), .C1(proc_wdata[19]), .Y(n3681) );
  AOI222X4 U265 ( .A0(mem_rdata[50]), .A1(n397), .B0(n3756), .B1(N137), .C0(
        n3757), .C1(proc_wdata[18]), .Y(n3682) );
  AOI222X4 U266 ( .A0(mem_rdata[49]), .A1(n398), .B0(n3756), .B1(N138), .C0(
        n3757), .C1(proc_wdata[17]), .Y(n3683) );
  AOI222X4 U267 ( .A0(mem_rdata[48]), .A1(n398), .B0(n3756), .B1(N139), .C0(
        n3757), .C1(proc_wdata[16]), .Y(n3684) );
  AOI222X4 U268 ( .A0(mem_rdata[47]), .A1(n397), .B0(n3756), .B1(N140), .C0(
        n3757), .C1(proc_wdata[15]), .Y(n3685) );
  AOI222X4 U269 ( .A0(mem_rdata[46]), .A1(n398), .B0(n3756), .B1(N141), .C0(
        n3757), .C1(proc_wdata[14]), .Y(n3686) );
  AOI222X4 U270 ( .A0(mem_rdata[45]), .A1(n398), .B0(n3756), .B1(N142), .C0(
        n3757), .C1(proc_wdata[13]), .Y(n3687) );
  AOI222X4 U271 ( .A0(mem_rdata[44]), .A1(n397), .B0(n3756), .B1(N143), .C0(
        n3757), .C1(proc_wdata[12]), .Y(n3688) );
  AOI222X4 U272 ( .A0(mem_rdata[43]), .A1(n397), .B0(n3756), .B1(N144), .C0(
        n3757), .C1(proc_wdata[11]), .Y(n3689) );
  AOI222X4 U273 ( .A0(mem_rdata[42]), .A1(n397), .B0(n3756), .B1(N145), .C0(
        n3757), .C1(proc_wdata[10]), .Y(n3690) );
  AOI222X4 U274 ( .A0(mem_rdata[41]), .A1(n397), .B0(n3756), .B1(N146), .C0(
        n3757), .C1(proc_wdata[9]), .Y(n3691) );
  AOI222X4 U275 ( .A0(mem_rdata[40]), .A1(n399), .B0(n3756), .B1(N147), .C0(
        n3757), .C1(proc_wdata[8]), .Y(n3692) );
  AOI222X4 U276 ( .A0(mem_rdata[39]), .A1(n399), .B0(n3756), .B1(N148), .C0(
        n3757), .C1(proc_wdata[7]), .Y(n3693) );
  AOI222X4 U277 ( .A0(mem_rdata[38]), .A1(n397), .B0(n3756), .B1(N149), .C0(
        n3757), .C1(proc_wdata[6]), .Y(n3694) );
  AOI222X4 U278 ( .A0(mem_rdata[37]), .A1(n399), .B0(n3756), .B1(N150), .C0(
        n3757), .C1(proc_wdata[5]), .Y(n3695) );
  AOI222X4 U279 ( .A0(mem_rdata[36]), .A1(n399), .B0(n3756), .B1(N151), .C0(
        n3757), .C1(proc_wdata[4]), .Y(n3696) );
  AOI222X4 U280 ( .A0(mem_rdata[35]), .A1(n397), .B0(n3756), .B1(N152), .C0(
        n3757), .C1(proc_wdata[3]), .Y(n3697) );
  AOI222X4 U281 ( .A0(mem_rdata[34]), .A1(n398), .B0(n3756), .B1(N153), .C0(
        n3757), .C1(proc_wdata[2]), .Y(n3698) );
  AOI222X4 U282 ( .A0(mem_rdata[33]), .A1(n399), .B0(n3756), .B1(N154), .C0(
        n3757), .C1(proc_wdata[1]), .Y(n3699) );
  AOI222X4 U283 ( .A0(mem_rdata[32]), .A1(n397), .B0(n3756), .B1(N155), .C0(
        n3757), .C1(proc_wdata[0]), .Y(n3700) );
  AOI222X4 U284 ( .A0(mem_rdata[31]), .A1(n399), .B0(n3759), .B1(N156), .C0(
        n3760), .C1(proc_wdata[31]), .Y(n3701) );
  AOI222X4 U285 ( .A0(mem_rdata[30]), .A1(n399), .B0(n3759), .B1(N157), .C0(
        n3760), .C1(proc_wdata[30]), .Y(n3702) );
  AOI222X4 U286 ( .A0(mem_rdata[29]), .A1(n397), .B0(n3759), .B1(N158), .C0(
        n3760), .C1(proc_wdata[29]), .Y(n3703) );
  AOI222X4 U287 ( .A0(mem_rdata[28]), .A1(n399), .B0(n3759), .B1(N159), .C0(
        n3760), .C1(proc_wdata[28]), .Y(n3704) );
  AOI222X4 U288 ( .A0(mem_rdata[27]), .A1(n399), .B0(n3759), .B1(N160), .C0(
        n3760), .C1(proc_wdata[27]), .Y(n3705) );
  AOI222X4 U289 ( .A0(mem_rdata[26]), .A1(n397), .B0(n3759), .B1(N161), .C0(
        n3760), .C1(proc_wdata[26]), .Y(n3706) );
  AOI222X4 U290 ( .A0(mem_rdata[25]), .A1(n400), .B0(n3759), .B1(N162), .C0(
        n3760), .C1(proc_wdata[25]), .Y(n3707) );
  AOI222X4 U291 ( .A0(mem_rdata[24]), .A1(n400), .B0(n3759), .B1(N163), .C0(
        n3760), .C1(proc_wdata[24]), .Y(n3708) );
  AOI222X4 U292 ( .A0(mem_rdata[23]), .A1(n398), .B0(n3759), .B1(N164), .C0(
        n3760), .C1(proc_wdata[23]), .Y(n3709) );
  AOI222X4 U293 ( .A0(mem_rdata[22]), .A1(n400), .B0(n3759), .B1(N165), .C0(
        n3760), .C1(proc_wdata[22]), .Y(n3710) );
  AOI222X4 U294 ( .A0(mem_rdata[21]), .A1(n400), .B0(n3759), .B1(N166), .C0(
        n3760), .C1(proc_wdata[21]), .Y(n3711) );
  AOI222X4 U295 ( .A0(mem_rdata[20]), .A1(n397), .B0(n3759), .B1(N167), .C0(
        n3760), .C1(proc_wdata[20]), .Y(n3712) );
  AOI222X4 U296 ( .A0(mem_rdata[19]), .A1(n400), .B0(n3759), .B1(N168), .C0(
        n3760), .C1(proc_wdata[19]), .Y(n3713) );
  AOI222X4 U297 ( .A0(mem_rdata[18]), .A1(n399), .B0(n3759), .B1(N169), .C0(
        n3760), .C1(proc_wdata[18]), .Y(n3714) );
  AOI222X4 U298 ( .A0(mem_rdata[17]), .A1(n398), .B0(n3759), .B1(N170), .C0(
        n3760), .C1(proc_wdata[17]), .Y(n3715) );
  AOI222X4 U299 ( .A0(mem_rdata[16]), .A1(n400), .B0(n3759), .B1(N171), .C0(
        n3760), .C1(proc_wdata[16]), .Y(n3716) );
  AOI222X4 U300 ( .A0(mem_rdata[15]), .A1(n400), .B0(n3759), .B1(N172), .C0(
        n3760), .C1(proc_wdata[15]), .Y(n3717) );
  AOI222X4 U301 ( .A0(mem_rdata[14]), .A1(n398), .B0(n3759), .B1(N173), .C0(
        n3760), .C1(proc_wdata[14]), .Y(n3718) );
  AOI222X4 U302 ( .A0(mem_rdata[13]), .A1(n400), .B0(n3759), .B1(N174), .C0(
        n3760), .C1(proc_wdata[13]), .Y(n3719) );
  AOI222X4 U303 ( .A0(mem_rdata[12]), .A1(n400), .B0(n3759), .B1(N175), .C0(
        n3760), .C1(proc_wdata[12]), .Y(n3720) );
  AOI222X4 U304 ( .A0(mem_rdata[11]), .A1(n398), .B0(n3759), .B1(N176), .C0(
        n3760), .C1(proc_wdata[11]), .Y(n3721) );
  AOI222X4 U305 ( .A0(mem_rdata[10]), .A1(n399), .B0(n3759), .B1(N177), .C0(
        n3760), .C1(proc_wdata[10]), .Y(n3722) );
  AOI222X4 U306 ( .A0(mem_rdata[9]), .A1(n400), .B0(n3759), .B1(N178), .C0(
        n3760), .C1(proc_wdata[9]), .Y(n3723) );
  AOI222X4 U307 ( .A0(mem_rdata[8]), .A1(n399), .B0(n3759), .B1(N179), .C0(
        n3760), .C1(proc_wdata[8]), .Y(n3724) );
  AOI222X4 U308 ( .A0(mem_rdata[7]), .A1(n400), .B0(n3759), .B1(N180), .C0(
        n3760), .C1(proc_wdata[7]), .Y(n3725) );
  AOI222X4 U309 ( .A0(mem_rdata[6]), .A1(n400), .B0(n3759), .B1(N181), .C0(
        n3760), .C1(proc_wdata[6]), .Y(n3726) );
  AOI222X4 U310 ( .A0(mem_rdata[5]), .A1(n399), .B0(n3759), .B1(N182), .C0(
        n3760), .C1(proc_wdata[5]), .Y(n3727) );
  AOI222X4 U311 ( .A0(mem_rdata[4]), .A1(n400), .B0(n3759), .B1(N183), .C0(
        n3760), .C1(proc_wdata[4]), .Y(n3728) );
  AOI222X4 U312 ( .A0(mem_rdata[3]), .A1(n400), .B0(n3759), .B1(N184), .C0(
        n3760), .C1(proc_wdata[3]), .Y(n3729) );
  AOI222X4 U313 ( .A0(mem_rdata[2]), .A1(n399), .B0(n3759), .B1(N185), .C0(
        n3760), .C1(proc_wdata[2]), .Y(n3730) );
  AOI222X4 U314 ( .A0(mem_rdata[1]), .A1(n3744), .B0(n3759), .B1(N186), .C0(
        n3760), .C1(proc_wdata[1]), .Y(n3731) );
  AOI222X4 U315 ( .A0(mem_rdata[0]), .A1(n396), .B0(n3759), .B1(N187), .C0(
        n3760), .C1(proc_wdata[0]), .Y(n3732) );
  INVX12 U316 ( .A(n8), .Y(mem_addr[9]) );
  INVX12 U317 ( .A(n7), .Y(mem_addr[8]) );
  INVX12 U318 ( .A(n6), .Y(mem_addr[7]) );
  INVX12 U319 ( .A(n5), .Y(mem_addr[6]) );
  INVX12 U320 ( .A(n4), .Y(mem_addr[5]) );
  INVX12 U321 ( .A(n3), .Y(mem_addr[4]) );
  INVX12 U322 ( .A(n2), .Y(mem_addr[3]) );
  INVX12 U323 ( .A(n26), .Y(mem_addr[27]) );
  INVX12 U324 ( .A(n25), .Y(mem_addr[26]) );
  INVX12 U325 ( .A(n24), .Y(mem_addr[25]) );
  INVX12 U326 ( .A(n23), .Y(mem_addr[24]) );
  INVX12 U327 ( .A(n22), .Y(mem_addr[23]) );
  INVX12 U328 ( .A(n21), .Y(mem_addr[22]) );
  INVX12 U329 ( .A(n20), .Y(mem_addr[21]) );
  INVX12 U330 ( .A(n19), .Y(mem_addr[20]) );
  INVX12 U331 ( .A(n18), .Y(mem_addr[19]) );
  INVX12 U332 ( .A(n17), .Y(mem_addr[18]) );
  INVX12 U333 ( .A(n16), .Y(mem_addr[17]) );
  INVX12 U334 ( .A(n15), .Y(mem_addr[16]) );
  INVX12 U335 ( .A(n14), .Y(mem_addr[15]) );
  INVX12 U336 ( .A(n13), .Y(mem_addr[14]) );
  INVX12 U337 ( .A(n12), .Y(mem_addr[13]) );
  INVX12 U338 ( .A(n11), .Y(mem_addr[12]) );
  INVX12 U339 ( .A(n10), .Y(mem_addr[11]) );
  INVX12 U340 ( .A(n9), .Y(mem_addr[10]) );
  INVX12 U341 ( .A(n36), .Y(mem_wdata[9]) );
  INVX12 U342 ( .A(n126), .Y(mem_wdata[99]) );
  INVX12 U343 ( .A(n125), .Y(mem_wdata[98]) );
  INVX12 U344 ( .A(n124), .Y(mem_wdata[97]) );
  INVX12 U345 ( .A(n123), .Y(mem_wdata[96]) );
  INVX12 U346 ( .A(n122), .Y(mem_wdata[95]) );
  INVX12 U347 ( .A(n121), .Y(mem_wdata[94]) );
  INVX12 U348 ( .A(n120), .Y(mem_wdata[93]) );
  INVX12 U349 ( .A(n119), .Y(mem_wdata[92]) );
  INVX12 U350 ( .A(n118), .Y(mem_wdata[91]) );
  INVX12 U351 ( .A(n117), .Y(mem_wdata[90]) );
  INVX12 U352 ( .A(n35), .Y(mem_wdata[8]) );
  INVX12 U353 ( .A(n116), .Y(mem_wdata[89]) );
  INVX12 U354 ( .A(n115), .Y(mem_wdata[88]) );
  INVX12 U355 ( .A(n114), .Y(mem_wdata[87]) );
  INVX12 U356 ( .A(n113), .Y(mem_wdata[86]) );
  INVX12 U357 ( .A(n112), .Y(mem_wdata[85]) );
  INVX12 U358 ( .A(n111), .Y(mem_wdata[84]) );
  INVX12 U359 ( .A(n110), .Y(mem_wdata[83]) );
  INVX12 U360 ( .A(n109), .Y(mem_wdata[82]) );
  INVX12 U361 ( .A(n108), .Y(mem_wdata[81]) );
  INVX12 U362 ( .A(n107), .Y(mem_wdata[80]) );
  INVX12 U363 ( .A(n34), .Y(mem_wdata[7]) );
  INVX12 U364 ( .A(n106), .Y(mem_wdata[79]) );
  INVX12 U365 ( .A(n105), .Y(mem_wdata[78]) );
  INVX12 U366 ( .A(n104), .Y(mem_wdata[77]) );
  INVX12 U367 ( .A(n103), .Y(mem_wdata[76]) );
  INVX12 U368 ( .A(n102), .Y(mem_wdata[75]) );
  INVX12 U369 ( .A(n101), .Y(mem_wdata[74]) );
  INVX12 U370 ( .A(n100), .Y(mem_wdata[73]) );
  INVX12 U371 ( .A(n99), .Y(mem_wdata[72]) );
  INVX12 U372 ( .A(n98), .Y(mem_wdata[71]) );
  INVX12 U373 ( .A(n97), .Y(mem_wdata[70]) );
  INVX12 U374 ( .A(n33), .Y(mem_wdata[6]) );
  INVX12 U375 ( .A(n96), .Y(mem_wdata[69]) );
  INVX12 U376 ( .A(n95), .Y(mem_wdata[68]) );
  INVX12 U377 ( .A(n94), .Y(mem_wdata[67]) );
  INVX12 U378 ( .A(n93), .Y(mem_wdata[66]) );
  INVX12 U379 ( .A(n92), .Y(mem_wdata[65]) );
  INVX12 U380 ( .A(n91), .Y(mem_wdata[64]) );
  INVX12 U381 ( .A(n90), .Y(mem_wdata[63]) );
  INVX12 U382 ( .A(n89), .Y(mem_wdata[62]) );
  INVX12 U383 ( .A(n88), .Y(mem_wdata[61]) );
  INVX12 U384 ( .A(n87), .Y(mem_wdata[60]) );
  INVX12 U385 ( .A(n32), .Y(mem_wdata[5]) );
  INVX12 U386 ( .A(n86), .Y(mem_wdata[59]) );
  INVX12 U387 ( .A(n85), .Y(mem_wdata[58]) );
  INVX12 U388 ( .A(n84), .Y(mem_wdata[57]) );
  INVX12 U389 ( .A(n83), .Y(mem_wdata[56]) );
  INVX12 U390 ( .A(n82), .Y(mem_wdata[55]) );
  INVX12 U391 ( .A(n81), .Y(mem_wdata[54]) );
  INVX12 U392 ( .A(n80), .Y(mem_wdata[53]) );
  INVX12 U393 ( .A(n79), .Y(mem_wdata[52]) );
  INVX12 U394 ( .A(n78), .Y(mem_wdata[51]) );
  INVX12 U395 ( .A(n77), .Y(mem_wdata[50]) );
  INVX12 U396 ( .A(n31), .Y(mem_wdata[4]) );
  INVX12 U397 ( .A(n76), .Y(mem_wdata[49]) );
  INVX12 U398 ( .A(n75), .Y(mem_wdata[48]) );
  INVX12 U399 ( .A(n74), .Y(mem_wdata[47]) );
  INVX12 U400 ( .A(n73), .Y(mem_wdata[46]) );
  INVX12 U401 ( .A(n72), .Y(mem_wdata[45]) );
  INVX12 U402 ( .A(n71), .Y(mem_wdata[44]) );
  INVX12 U403 ( .A(n70), .Y(mem_wdata[43]) );
  INVX12 U404 ( .A(n69), .Y(mem_wdata[42]) );
  INVX12 U405 ( .A(n68), .Y(mem_wdata[41]) );
  INVX12 U406 ( .A(n67), .Y(mem_wdata[40]) );
  INVX12 U407 ( .A(n30), .Y(mem_wdata[3]) );
  INVX12 U408 ( .A(n66), .Y(mem_wdata[39]) );
  INVX12 U409 ( .A(n65), .Y(mem_wdata[38]) );
  INVX12 U410 ( .A(n64), .Y(mem_wdata[37]) );
  INVX12 U411 ( .A(n63), .Y(mem_wdata[36]) );
  INVX12 U412 ( .A(n62), .Y(mem_wdata[35]) );
  INVX12 U413 ( .A(n61), .Y(mem_wdata[34]) );
  INVX12 U414 ( .A(n60), .Y(mem_wdata[33]) );
  INVX12 U415 ( .A(n59), .Y(mem_wdata[32]) );
  INVX12 U416 ( .A(n58), .Y(mem_wdata[31]) );
  INVX12 U417 ( .A(n57), .Y(mem_wdata[30]) );
  INVX12 U418 ( .A(n29), .Y(mem_wdata[2]) );
  INVX12 U419 ( .A(n56), .Y(mem_wdata[29]) );
  INVX12 U420 ( .A(n55), .Y(mem_wdata[28]) );
  INVX12 U421 ( .A(n54), .Y(mem_wdata[27]) );
  INVX12 U422 ( .A(n53), .Y(mem_wdata[26]) );
  INVX12 U423 ( .A(n52), .Y(mem_wdata[25]) );
  INVX12 U424 ( .A(n51), .Y(mem_wdata[24]) );
  INVX12 U425 ( .A(n50), .Y(mem_wdata[23]) );
  INVX12 U426 ( .A(n49), .Y(mem_wdata[22]) );
  INVX12 U427 ( .A(n48), .Y(mem_wdata[21]) );
  INVX12 U428 ( .A(n47), .Y(mem_wdata[20]) );
  INVX12 U429 ( .A(n28), .Y(mem_wdata[1]) );
  INVX12 U430 ( .A(n46), .Y(mem_wdata[19]) );
  INVX12 U431 ( .A(n45), .Y(mem_wdata[18]) );
  INVX12 U432 ( .A(n44), .Y(mem_wdata[17]) );
  INVX12 U433 ( .A(n43), .Y(mem_wdata[16]) );
  INVX12 U434 ( .A(n42), .Y(mem_wdata[15]) );
  INVX12 U435 ( .A(n41), .Y(mem_wdata[14]) );
  INVX12 U436 ( .A(n40), .Y(mem_wdata[13]) );
  INVX12 U437 ( .A(n39), .Y(mem_wdata[12]) );
  INVX12 U438 ( .A(n154), .Y(mem_wdata[127]) );
  INVX12 U439 ( .A(n153), .Y(mem_wdata[126]) );
  INVX12 U440 ( .A(n152), .Y(mem_wdata[125]) );
  INVX12 U441 ( .A(n151), .Y(mem_wdata[124]) );
  INVX12 U442 ( .A(n150), .Y(mem_wdata[123]) );
  INVX12 U443 ( .A(n149), .Y(mem_wdata[122]) );
  INVX12 U444 ( .A(n148), .Y(mem_wdata[121]) );
  INVX12 U445 ( .A(n147), .Y(mem_wdata[120]) );
  INVX12 U446 ( .A(n38), .Y(mem_wdata[11]) );
  INVX12 U447 ( .A(n146), .Y(mem_wdata[119]) );
  INVX12 U448 ( .A(n145), .Y(mem_wdata[118]) );
  INVX12 U449 ( .A(n144), .Y(mem_wdata[117]) );
  INVX12 U450 ( .A(n143), .Y(mem_wdata[116]) );
  INVX12 U451 ( .A(n142), .Y(mem_wdata[115]) );
  INVX12 U452 ( .A(n141), .Y(mem_wdata[114]) );
  INVX12 U453 ( .A(n140), .Y(mem_wdata[113]) );
  INVX12 U454 ( .A(n139), .Y(mem_wdata[112]) );
  INVX12 U455 ( .A(n138), .Y(mem_wdata[111]) );
  INVX12 U456 ( .A(n137), .Y(mem_wdata[110]) );
  INVX12 U457 ( .A(n37), .Y(mem_wdata[10]) );
  INVX12 U458 ( .A(n136), .Y(mem_wdata[109]) );
  INVX12 U459 ( .A(n135), .Y(mem_wdata[108]) );
  INVX12 U460 ( .A(n134), .Y(mem_wdata[107]) );
  INVX12 U461 ( .A(n133), .Y(mem_wdata[106]) );
  INVX12 U462 ( .A(n132), .Y(mem_wdata[105]) );
  INVX12 U463 ( .A(n131), .Y(mem_wdata[104]) );
  INVX12 U464 ( .A(n130), .Y(mem_wdata[103]) );
  INVX12 U465 ( .A(n129), .Y(mem_wdata[102]) );
  INVX12 U466 ( .A(n128), .Y(mem_wdata[101]) );
  INVX12 U467 ( .A(n127), .Y(mem_wdata[100]) );
  INVX12 U468 ( .A(n27), .Y(mem_wdata[0]) );
  INVX12 U469 ( .A(n1), .Y(mem_addr[2]) );
  INVX12 U470 ( .A(n156), .Y(mem_addr[1]) );
  INVX12 U471 ( .A(n155), .Y(mem_addr[0]) );
  NAND3X6 U472 ( .A(proc_addr[0]), .B(n3574), .C(proc_addr[1]), .Y(n3417) );
  BUFX4 U473 ( .A(n3745), .Y(n316) );
  AOI22X2 U474 ( .A0(proc_addr[8]), .A1(n398), .B0(n3745), .B1(N56), .Y(n3601)
         );
  AOI22X2 U475 ( .A0(proc_addr[9]), .A1(n396), .B0(n3745), .B1(N55), .Y(n3600)
         );
  AOI22X2 U476 ( .A0(proc_addr[10]), .A1(n399), .B0(n3745), .B1(N54), .Y(n3599) );
  NOR3X6 U477 ( .A(n3576), .B(n3575), .C(n3742), .Y(n3749) );
  CLKINVX1 U478 ( .A(n3804), .Y(n317) );
  INVX16 U479 ( .A(n317), .Y(mem_read) );
  NAND2X6 U480 ( .A(proc_addr[1]), .B(n158), .Y(n3411) );
  INVX3 U481 ( .A(proc_addr[0]), .Y(n3575) );
  NAND2X6 U482 ( .A(proc_addr[0]), .B(n159), .Y(n3413) );
  INVX3 U483 ( .A(proc_addr[1]), .Y(n3576) );
  OAI221X1 U484 ( .A0(n3410), .A1(n3746), .B0(mem_ready), .B1(n3764), .C0(
        n3747), .Y(n3751) );
  INVX6 U485 ( .A(n3761), .Y(n3759) );
  INVX6 U486 ( .A(n3755), .Y(n3754) );
  INVX6 U487 ( .A(n3758), .Y(n3756) );
  INVX6 U488 ( .A(n3750), .Y(n3748) );
  NOR2X2 U489 ( .A(n3766), .B(n3763), .Y(n3574) );
  AOI211X4 U490 ( .A0(proc_read), .A1(mem_ready), .B0(n3740), .C0(N33), .Y(
        n3577) );
  CLKINVX2 U491 ( .A(n3740), .Y(n3742) );
  AND2X2 U492 ( .A(n3741), .B(n3742), .Y(n3579) );
  OA22XL U493 ( .A0(n157), .A1(n3572), .B0(n3417), .B1(n3573), .Y(n3571) );
  OA22XL U494 ( .A0(n157), .A1(n3517), .B0(n3417), .B1(n3518), .Y(n3516) );
  OA22XL U495 ( .A0(n157), .A1(n3462), .B0(n3417), .B1(n3463), .Y(n3461) );
  OA22XL U496 ( .A0(n157), .A1(n3447), .B0(n3417), .B1(n3448), .Y(n3446) );
  OA22XL U497 ( .A0(n157), .A1(n3442), .B0(n3417), .B1(n3443), .Y(n3441) );
  OA22XL U498 ( .A0(n157), .A1(n3437), .B0(n3417), .B1(n3438), .Y(n3436) );
  OA22XL U499 ( .A0(n157), .A1(n3432), .B0(n3417), .B1(n3433), .Y(n3431) );
  OA22XL U500 ( .A0(n157), .A1(n3427), .B0(n3417), .B1(n3428), .Y(n3426) );
  OA22XL U501 ( .A0(n157), .A1(n3422), .B0(n3417), .B1(n3423), .Y(n3421) );
  OA22XL U502 ( .A0(n157), .A1(n3416), .B0(n3417), .B1(n3418), .Y(n3415) );
  OA22XL U503 ( .A0(n157), .A1(n3567), .B0(n3417), .B1(n3568), .Y(n3566) );
  OA22XL U504 ( .A0(n157), .A1(n3562), .B0(n3417), .B1(n3563), .Y(n3561) );
  OA22XL U505 ( .A0(n157), .A1(n3557), .B0(n3417), .B1(n3558), .Y(n3556) );
  OA22XL U506 ( .A0(n157), .A1(n3552), .B0(n3417), .B1(n3553), .Y(n3551) );
  OA22XL U507 ( .A0(n157), .A1(n3547), .B0(n3417), .B1(n3548), .Y(n3546) );
  OA22XL U508 ( .A0(n157), .A1(n3542), .B0(n3417), .B1(n3543), .Y(n3541) );
  OA22XL U509 ( .A0(n157), .A1(n3537), .B0(n3417), .B1(n3538), .Y(n3536) );
  OA22XL U510 ( .A0(n157), .A1(n3532), .B0(n3417), .B1(n3533), .Y(n3531) );
  OA22XL U511 ( .A0(n157), .A1(n3527), .B0(n3417), .B1(n3528), .Y(n3526) );
  OA22XL U512 ( .A0(n157), .A1(n3522), .B0(n3417), .B1(n3523), .Y(n3521) );
  OA22XL U513 ( .A0(n157), .A1(n3512), .B0(n3417), .B1(n3513), .Y(n3511) );
  OA22XL U514 ( .A0(n157), .A1(n3507), .B0(n3417), .B1(n3508), .Y(n3506) );
  OA22XL U515 ( .A0(n157), .A1(n3502), .B0(n3417), .B1(n3503), .Y(n3501) );
  OA22XL U516 ( .A0(n157), .A1(n3497), .B0(n3417), .B1(n3498), .Y(n3496) );
  OA22XL U517 ( .A0(n157), .A1(n3492), .B0(n3417), .B1(n3493), .Y(n3491) );
  OA22XL U518 ( .A0(n157), .A1(n3487), .B0(n3417), .B1(n3488), .Y(n3486) );
  OA22XL U519 ( .A0(n157), .A1(n3482), .B0(n3417), .B1(n3483), .Y(n3481) );
  OA22XL U520 ( .A0(n157), .A1(n3477), .B0(n3417), .B1(n3478), .Y(n3476) );
  OA22XL U521 ( .A0(n157), .A1(n3472), .B0(n3417), .B1(n3473), .Y(n3471) );
  OA22XL U522 ( .A0(n157), .A1(n3467), .B0(n3417), .B1(n3468), .Y(n3466) );
  OA22XL U523 ( .A0(n157), .A1(n3457), .B0(n3417), .B1(n3458), .Y(n3456) );
  OA22XL U524 ( .A0(n157), .A1(n3452), .B0(n3417), .B1(n3453), .Y(n3451) );
  AOI211XL U525 ( .A0(n3765), .A1(N34), .B0(n3574), .C0(n3408), .Y(n3747) );
  XNOR2XL U526 ( .A(N38), .B(proc_addr[26]), .Y(n3779) );
  XNOR2XL U527 ( .A(N54), .B(proc_addr[10]), .Y(n3801) );
  XNOR2XL U528 ( .A(N56), .B(proc_addr[8]), .Y(n3802) );
  XNOR2XL U529 ( .A(N55), .B(proc_addr[9]), .Y(n3803) );
  MXI2XL U530 ( .A(n541), .B(n3732), .S0(n385), .Y(n1781) );
  MXI2XL U531 ( .A(n542), .B(n3731), .S0(n385), .Y(n1782) );
  MXI2XL U532 ( .A(n543), .B(n3730), .S0(n385), .Y(n1783) );
  MXI2XL U533 ( .A(n544), .B(n3729), .S0(n385), .Y(n1784) );
  MXI2XL U534 ( .A(n545), .B(n3728), .S0(n385), .Y(n1785) );
  MXI2XL U535 ( .A(n546), .B(n3727), .S0(n385), .Y(n1786) );
  MXI2XL U536 ( .A(n547), .B(n3726), .S0(n385), .Y(n1787) );
  MXI2XL U537 ( .A(n548), .B(n3725), .S0(n385), .Y(n1788) );
  MXI2XL U538 ( .A(n549), .B(n3724), .S0(n385), .Y(n1789) );
  MXI2XL U539 ( .A(n550), .B(n3723), .S0(n385), .Y(n1790) );
  MXI2XL U540 ( .A(n551), .B(n3722), .S0(n385), .Y(n1791) );
  MXI2XL U541 ( .A(n552), .B(n3721), .S0(n385), .Y(n1792) );
  MXI2XL U542 ( .A(n553), .B(n3720), .S0(n385), .Y(n1793) );
  MXI2XL U543 ( .A(n554), .B(n3719), .S0(n386), .Y(n1794) );
  MXI2XL U544 ( .A(n555), .B(n3718), .S0(n386), .Y(n1795) );
  MXI2XL U545 ( .A(n556), .B(n3717), .S0(n386), .Y(n1796) );
  MXI2XL U546 ( .A(n557), .B(n3716), .S0(n386), .Y(n1797) );
  MXI2XL U547 ( .A(n558), .B(n3715), .S0(n386), .Y(n1798) );
  MXI2XL U548 ( .A(n559), .B(n3714), .S0(n386), .Y(n1799) );
  MXI2XL U549 ( .A(n560), .B(n3713), .S0(n386), .Y(n1800) );
  MXI2XL U550 ( .A(n561), .B(n3712), .S0(n386), .Y(n1801) );
  MXI2XL U551 ( .A(n562), .B(n3711), .S0(n386), .Y(n1802) );
  MXI2XL U552 ( .A(n563), .B(n3710), .S0(n386), .Y(n1803) );
  MXI2XL U553 ( .A(n564), .B(n3709), .S0(n386), .Y(n1804) );
  MXI2XL U554 ( .A(n565), .B(n3708), .S0(n386), .Y(n1805) );
  MXI2XL U555 ( .A(n566), .B(n3707), .S0(n386), .Y(n1806) );
  MXI2XL U556 ( .A(n567), .B(n3706), .S0(n387), .Y(n1807) );
  MXI2XL U557 ( .A(n568), .B(n3705), .S0(n387), .Y(n1808) );
  MXI2XL U558 ( .A(n569), .B(n3704), .S0(n387), .Y(n1809) );
  MXI2XL U559 ( .A(n570), .B(n3703), .S0(n387), .Y(n1810) );
  MXI2XL U560 ( .A(n571), .B(n3702), .S0(n387), .Y(n1811) );
  MXI2XL U561 ( .A(n572), .B(n3701), .S0(n387), .Y(n1812) );
  MXI2XL U562 ( .A(n573), .B(n3700), .S0(n387), .Y(n1813) );
  MXI2XL U563 ( .A(n574), .B(n3699), .S0(n387), .Y(n1814) );
  MXI2XL U564 ( .A(n575), .B(n3698), .S0(n387), .Y(n1815) );
  MXI2XL U565 ( .A(n576), .B(n3697), .S0(n387), .Y(n1816) );
  MXI2XL U566 ( .A(n577), .B(n3696), .S0(n387), .Y(n1817) );
  MXI2XL U567 ( .A(n578), .B(n3695), .S0(n387), .Y(n1818) );
  MXI2XL U568 ( .A(n579), .B(n3694), .S0(n387), .Y(n1819) );
  MXI2XL U569 ( .A(n580), .B(n3693), .S0(n388), .Y(n1820) );
  MXI2XL U570 ( .A(n581), .B(n3692), .S0(n388), .Y(n1821) );
  MXI2XL U571 ( .A(n582), .B(n3691), .S0(n388), .Y(n1822) );
  MXI2XL U572 ( .A(n583), .B(n3690), .S0(n388), .Y(n1823) );
  MXI2XL U573 ( .A(n584), .B(n3689), .S0(n388), .Y(n1824) );
  MXI2XL U574 ( .A(n585), .B(n3688), .S0(n388), .Y(n1825) );
  MXI2XL U575 ( .A(n586), .B(n3687), .S0(n388), .Y(n1826) );
  MXI2XL U576 ( .A(n587), .B(n3686), .S0(n388), .Y(n1827) );
  MXI2XL U577 ( .A(n588), .B(n3685), .S0(n388), .Y(n1828) );
  MXI2XL U578 ( .A(n589), .B(n3684), .S0(n388), .Y(n1829) );
  MXI2XL U579 ( .A(n590), .B(n3683), .S0(n388), .Y(n1830) );
  MXI2XL U580 ( .A(n591), .B(n3682), .S0(n388), .Y(n1831) );
  MXI2XL U581 ( .A(n592), .B(n3681), .S0(n388), .Y(n1832) );
  MXI2XL U582 ( .A(n593), .B(n3680), .S0(n389), .Y(n1833) );
  MXI2XL U583 ( .A(n594), .B(n3679), .S0(n389), .Y(n1834) );
  MXI2XL U584 ( .A(n595), .B(n3678), .S0(n389), .Y(n1835) );
  MXI2XL U585 ( .A(n596), .B(n3677), .S0(n389), .Y(n1836) );
  MXI2XL U586 ( .A(n597), .B(n3676), .S0(n389), .Y(n1837) );
  MXI2XL U587 ( .A(n598), .B(n3675), .S0(n389), .Y(n1838) );
  MXI2XL U588 ( .A(n599), .B(n3674), .S0(n389), .Y(n1839) );
  MXI2XL U589 ( .A(n600), .B(n3673), .S0(n389), .Y(n1840) );
  MXI2XL U590 ( .A(n601), .B(n3672), .S0(n389), .Y(n1841) );
  MXI2XL U591 ( .A(n602), .B(n3671), .S0(n389), .Y(n1842) );
  MXI2XL U592 ( .A(n603), .B(n3670), .S0(n389), .Y(n1843) );
  MXI2XL U593 ( .A(n604), .B(n3669), .S0(n389), .Y(n1844) );
  MXI2XL U594 ( .A(n637), .B(n3636), .S0(n3739), .Y(n1877) );
  MXI2XL U595 ( .A(n638), .B(n3635), .S0(n387), .Y(n1878) );
  MXI2XL U596 ( .A(n639), .B(n3634), .S0(n391), .Y(n1879) );
  MXI2XL U597 ( .A(n640), .B(n3633), .S0(n388), .Y(n1880) );
  MXI2XL U598 ( .A(n641), .B(n3632), .S0(n392), .Y(n1881) );
  MXI2XL U599 ( .A(n642), .B(n3631), .S0(n385), .Y(n1882) );
  MXI2XL U600 ( .A(n643), .B(n3630), .S0(n386), .Y(n1883) );
  MXI2XL U601 ( .A(n644), .B(n3629), .S0(n389), .Y(n1884) );
  MXI2XL U602 ( .A(n645), .B(n3628), .S0(n392), .Y(n1885) );
  MXI2XL U603 ( .A(n646), .B(n3627), .S0(n392), .Y(n1886) );
  MXI2XL U604 ( .A(n647), .B(n3626), .S0(n392), .Y(n1887) );
  MXI2XL U605 ( .A(n648), .B(n3625), .S0(n392), .Y(n1888) );
  MXI2XL U606 ( .A(n649), .B(n3624), .S0(n392), .Y(n1889) );
  MXI2XL U607 ( .A(n650), .B(n3623), .S0(n392), .Y(n1890) );
  MXI2XL U608 ( .A(n651), .B(n3622), .S0(n392), .Y(n1891) );
  MXI2XL U609 ( .A(n652), .B(n3621), .S0(n392), .Y(n1892) );
  MXI2XL U610 ( .A(n653), .B(n3620), .S0(n392), .Y(n1893) );
  MXI2XL U611 ( .A(n654), .B(n3619), .S0(n392), .Y(n1894) );
  MXI2XL U612 ( .A(n655), .B(n3618), .S0(n392), .Y(n1895) );
  MXI2XL U613 ( .A(n656), .B(n3617), .S0(n392), .Y(n1896) );
  MXI2XL U614 ( .A(n657), .B(n3616), .S0(n392), .Y(n1897) );
  MXI2XL U615 ( .A(n658), .B(n3615), .S0(n386), .Y(n1898) );
  MXI2XL U616 ( .A(n659), .B(n3614), .S0(n389), .Y(n1899) );
  MXI2XL U617 ( .A(n660), .B(n3613), .S0(n393), .Y(n1900) );
  MXI2XL U618 ( .A(n661), .B(n3612), .S0(n3739), .Y(n1901) );
  MXI2XL U619 ( .A(n662), .B(n3611), .S0(n390), .Y(n1902) );
  MXI2XL U620 ( .A(n663), .B(n3610), .S0(n387), .Y(n1903) );
  MXI2XL U621 ( .A(n664), .B(n3609), .S0(n391), .Y(n1904) );
  MXI2XL U622 ( .A(n665), .B(n3608), .S0(n388), .Y(n1905) );
  MXI2XL U623 ( .A(n666), .B(n3607), .S0(n392), .Y(n1906) );
  MXI2XL U624 ( .A(n667), .B(n3606), .S0(n385), .Y(n1907) );
  MXI2XL U625 ( .A(n668), .B(n3605), .S0(n386), .Y(n1908) );
  MXI2XL U626 ( .A(n696), .B(n3732), .S0(n376), .Y(n1936) );
  MXI2XL U627 ( .A(n697), .B(n3731), .S0(n376), .Y(n1937) );
  MXI2XL U628 ( .A(n698), .B(n3730), .S0(n376), .Y(n1938) );
  MXI2XL U629 ( .A(n699), .B(n3729), .S0(n376), .Y(n1939) );
  MXI2XL U630 ( .A(n700), .B(n3728), .S0(n376), .Y(n1940) );
  MXI2XL U631 ( .A(n701), .B(n3727), .S0(n376), .Y(n1941) );
  MXI2XL U632 ( .A(n702), .B(n3726), .S0(n376), .Y(n1942) );
  MXI2XL U633 ( .A(n703), .B(n3725), .S0(n376), .Y(n1943) );
  MXI2XL U634 ( .A(n704), .B(n3724), .S0(n376), .Y(n1944) );
  MXI2XL U635 ( .A(n705), .B(n3723), .S0(n376), .Y(n1945) );
  MXI2XL U636 ( .A(n706), .B(n3722), .S0(n376), .Y(n1946) );
  MXI2XL U637 ( .A(n707), .B(n3721), .S0(n376), .Y(n1947) );
  MXI2XL U638 ( .A(n708), .B(n3720), .S0(n376), .Y(n1948) );
  MXI2XL U639 ( .A(n709), .B(n3719), .S0(n377), .Y(n1949) );
  MXI2XL U640 ( .A(n710), .B(n3718), .S0(n377), .Y(n1950) );
  MXI2XL U641 ( .A(n711), .B(n3717), .S0(n377), .Y(n1951) );
  MXI2XL U642 ( .A(n712), .B(n3716), .S0(n377), .Y(n1952) );
  MXI2XL U643 ( .A(n713), .B(n3715), .S0(n377), .Y(n1953) );
  MXI2XL U644 ( .A(n714), .B(n3714), .S0(n377), .Y(n1954) );
  MXI2XL U645 ( .A(n715), .B(n3713), .S0(n377), .Y(n1955) );
  MXI2XL U646 ( .A(n716), .B(n3712), .S0(n377), .Y(n1956) );
  MXI2XL U647 ( .A(n717), .B(n3711), .S0(n377), .Y(n1957) );
  MXI2XL U648 ( .A(n718), .B(n3710), .S0(n377), .Y(n1958) );
  MXI2XL U649 ( .A(n719), .B(n3709), .S0(n377), .Y(n1959) );
  MXI2XL U650 ( .A(n720), .B(n3708), .S0(n377), .Y(n1960) );
  MXI2XL U651 ( .A(n721), .B(n3707), .S0(n377), .Y(n1961) );
  MXI2XL U652 ( .A(n722), .B(n3706), .S0(n378), .Y(n1962) );
  MXI2XL U653 ( .A(n723), .B(n3705), .S0(n378), .Y(n1963) );
  MXI2XL U654 ( .A(n724), .B(n3704), .S0(n378), .Y(n1964) );
  MXI2XL U655 ( .A(n725), .B(n3703), .S0(n378), .Y(n1965) );
  MXI2XL U656 ( .A(n726), .B(n3702), .S0(n378), .Y(n1966) );
  MXI2XL U657 ( .A(n727), .B(n3701), .S0(n378), .Y(n1967) );
  MXI2XL U658 ( .A(n728), .B(n3700), .S0(n378), .Y(n1968) );
  MXI2XL U659 ( .A(n729), .B(n3699), .S0(n378), .Y(n1969) );
  MXI2XL U660 ( .A(n730), .B(n3698), .S0(n378), .Y(n1970) );
  MXI2XL U661 ( .A(n731), .B(n3697), .S0(n378), .Y(n1971) );
  MXI2XL U662 ( .A(n732), .B(n3696), .S0(n378), .Y(n1972) );
  MXI2XL U663 ( .A(n733), .B(n3695), .S0(n378), .Y(n1973) );
  MXI2XL U664 ( .A(n734), .B(n3694), .S0(n378), .Y(n1974) );
  MXI2XL U665 ( .A(n735), .B(n3693), .S0(n379), .Y(n1975) );
  MXI2XL U666 ( .A(n736), .B(n3692), .S0(n379), .Y(n1976) );
  MXI2XL U667 ( .A(n737), .B(n3691), .S0(n379), .Y(n1977) );
  MXI2XL U668 ( .A(n738), .B(n3690), .S0(n379), .Y(n1978) );
  MXI2XL U669 ( .A(n739), .B(n3689), .S0(n379), .Y(n1979) );
  MXI2XL U670 ( .A(n740), .B(n3688), .S0(n379), .Y(n1980) );
  MXI2XL U671 ( .A(n741), .B(n3687), .S0(n379), .Y(n1981) );
  MXI2XL U672 ( .A(n742), .B(n3686), .S0(n379), .Y(n1982) );
  MXI2XL U673 ( .A(n743), .B(n3685), .S0(n379), .Y(n1983) );
  MXI2XL U674 ( .A(n744), .B(n3684), .S0(n379), .Y(n1984) );
  MXI2XL U675 ( .A(n745), .B(n3683), .S0(n379), .Y(n1985) );
  MXI2XL U676 ( .A(n746), .B(n3682), .S0(n379), .Y(n1986) );
  MXI2XL U677 ( .A(n747), .B(n3681), .S0(n379), .Y(n1987) );
  MXI2XL U678 ( .A(n748), .B(n3680), .S0(n380), .Y(n1988) );
  MXI2XL U679 ( .A(n749), .B(n3679), .S0(n380), .Y(n1989) );
  MXI2XL U680 ( .A(n750), .B(n3678), .S0(n380), .Y(n1990) );
  MXI2XL U681 ( .A(n751), .B(n3677), .S0(n380), .Y(n1991) );
  MXI2XL U682 ( .A(n752), .B(n3676), .S0(n380), .Y(n1992) );
  MXI2XL U683 ( .A(n753), .B(n3675), .S0(n380), .Y(n1993) );
  MXI2XL U684 ( .A(n754), .B(n3674), .S0(n380), .Y(n1994) );
  MXI2XL U685 ( .A(n755), .B(n3673), .S0(n380), .Y(n1995) );
  MXI2XL U686 ( .A(n756), .B(n3672), .S0(n380), .Y(n1996) );
  MXI2XL U687 ( .A(n757), .B(n3671), .S0(n380), .Y(n1997) );
  MXI2XL U688 ( .A(n758), .B(n3670), .S0(n380), .Y(n1998) );
  MXI2XL U689 ( .A(n759), .B(n3669), .S0(n380), .Y(n1999) );
  MXI2XL U690 ( .A(n792), .B(n3636), .S0(n3738), .Y(n2032) );
  MXI2XL U691 ( .A(n793), .B(n3635), .S0(n378), .Y(n2033) );
  MXI2XL U692 ( .A(n794), .B(n3634), .S0(n382), .Y(n2034) );
  MXI2XL U693 ( .A(n795), .B(n3633), .S0(n379), .Y(n2035) );
  MXI2XL U694 ( .A(n796), .B(n3632), .S0(n383), .Y(n2036) );
  MXI2XL U695 ( .A(n797), .B(n3631), .S0(n376), .Y(n2037) );
  MXI2XL U696 ( .A(n798), .B(n3630), .S0(n377), .Y(n2038) );
  MXI2XL U697 ( .A(n799), .B(n3629), .S0(n380), .Y(n2039) );
  MXI2XL U698 ( .A(n800), .B(n3628), .S0(n383), .Y(n2040) );
  MXI2XL U699 ( .A(n801), .B(n3627), .S0(n383), .Y(n2041) );
  MXI2XL U700 ( .A(n802), .B(n3626), .S0(n383), .Y(n2042) );
  MXI2XL U701 ( .A(n803), .B(n3625), .S0(n383), .Y(n2043) );
  MXI2XL U702 ( .A(n804), .B(n3624), .S0(n383), .Y(n2044) );
  MXI2XL U703 ( .A(n805), .B(n3623), .S0(n383), .Y(n2045) );
  MXI2XL U704 ( .A(n806), .B(n3622), .S0(n383), .Y(n2046) );
  MXI2XL U705 ( .A(n807), .B(n3621), .S0(n383), .Y(n2047) );
  MXI2XL U706 ( .A(n808), .B(n3620), .S0(n383), .Y(n2048) );
  MXI2XL U707 ( .A(n809), .B(n3619), .S0(n383), .Y(n2049) );
  MXI2XL U708 ( .A(n810), .B(n3618), .S0(n383), .Y(n2050) );
  MXI2XL U709 ( .A(n811), .B(n3617), .S0(n383), .Y(n2051) );
  MXI2XL U710 ( .A(n812), .B(n3616), .S0(n383), .Y(n2052) );
  MXI2XL U711 ( .A(n813), .B(n3615), .S0(n377), .Y(n2053) );
  MXI2XL U712 ( .A(n814), .B(n3614), .S0(n380), .Y(n2054) );
  MXI2XL U713 ( .A(n815), .B(n3613), .S0(n384), .Y(n2055) );
  MXI2XL U714 ( .A(n816), .B(n3612), .S0(n3738), .Y(n2056) );
  MXI2XL U715 ( .A(n817), .B(n3611), .S0(n381), .Y(n2057) );
  MXI2XL U716 ( .A(n818), .B(n3610), .S0(n378), .Y(n2058) );
  MXI2XL U717 ( .A(n819), .B(n3609), .S0(n382), .Y(n2059) );
  MXI2XL U718 ( .A(n820), .B(n3608), .S0(n379), .Y(n2060) );
  MXI2XL U719 ( .A(n821), .B(n3607), .S0(n383), .Y(n2061) );
  MXI2XL U720 ( .A(n822), .B(n3606), .S0(n376), .Y(n2062) );
  MXI2XL U721 ( .A(n823), .B(n3605), .S0(n377), .Y(n2063) );
  MXI2XL U722 ( .A(n851), .B(n3732), .S0(n367), .Y(n2091) );
  MXI2XL U723 ( .A(n852), .B(n3731), .S0(n367), .Y(n2092) );
  MXI2XL U724 ( .A(n853), .B(n3730), .S0(n367), .Y(n2093) );
  MXI2XL U725 ( .A(n854), .B(n3729), .S0(n367), .Y(n2094) );
  MXI2XL U726 ( .A(n855), .B(n3728), .S0(n367), .Y(n2095) );
  MXI2XL U727 ( .A(n856), .B(n3727), .S0(n367), .Y(n2096) );
  MXI2XL U728 ( .A(n857), .B(n3726), .S0(n367), .Y(n2097) );
  MXI2XL U729 ( .A(n858), .B(n3725), .S0(n367), .Y(n2098) );
  MXI2XL U730 ( .A(n859), .B(n3724), .S0(n367), .Y(n2099) );
  MXI2XL U731 ( .A(n860), .B(n3723), .S0(n367), .Y(n2100) );
  MXI2XL U732 ( .A(n861), .B(n3722), .S0(n367), .Y(n2101) );
  MXI2XL U733 ( .A(n862), .B(n3721), .S0(n367), .Y(n2102) );
  MXI2XL U734 ( .A(n863), .B(n3720), .S0(n367), .Y(n2103) );
  MXI2XL U735 ( .A(n864), .B(n3719), .S0(n368), .Y(n2104) );
  MXI2XL U736 ( .A(n865), .B(n3718), .S0(n368), .Y(n2105) );
  MXI2XL U737 ( .A(n866), .B(n3717), .S0(n368), .Y(n2106) );
  MXI2XL U738 ( .A(n867), .B(n3716), .S0(n368), .Y(n2107) );
  MXI2XL U739 ( .A(n868), .B(n3715), .S0(n368), .Y(n2108) );
  MXI2XL U740 ( .A(n869), .B(n3714), .S0(n368), .Y(n2109) );
  MXI2XL U741 ( .A(n870), .B(n3713), .S0(n368), .Y(n2110) );
  MXI2XL U742 ( .A(n871), .B(n3712), .S0(n368), .Y(n2111) );
  MXI2XL U743 ( .A(n872), .B(n3711), .S0(n368), .Y(n2112) );
  MXI2XL U744 ( .A(n873), .B(n3710), .S0(n368), .Y(n2113) );
  MXI2XL U745 ( .A(n874), .B(n3709), .S0(n368), .Y(n2114) );
  MXI2XL U746 ( .A(n875), .B(n3708), .S0(n368), .Y(n2115) );
  MXI2XL U747 ( .A(n876), .B(n3707), .S0(n368), .Y(n2116) );
  MXI2XL U748 ( .A(n877), .B(n3706), .S0(n369), .Y(n2117) );
  MXI2XL U749 ( .A(n878), .B(n3705), .S0(n369), .Y(n2118) );
  MXI2XL U750 ( .A(n879), .B(n3704), .S0(n369), .Y(n2119) );
  MXI2XL U751 ( .A(n880), .B(n3703), .S0(n369), .Y(n2120) );
  MXI2XL U752 ( .A(n881), .B(n3702), .S0(n369), .Y(n2121) );
  MXI2XL U753 ( .A(n882), .B(n3701), .S0(n369), .Y(n2122) );
  MXI2XL U754 ( .A(n883), .B(n3700), .S0(n369), .Y(n2123) );
  MXI2XL U755 ( .A(n884), .B(n3699), .S0(n369), .Y(n2124) );
  MXI2XL U756 ( .A(n885), .B(n3698), .S0(n369), .Y(n2125) );
  MXI2XL U757 ( .A(n886), .B(n3697), .S0(n369), .Y(n2126) );
  MXI2XL U758 ( .A(n887), .B(n3696), .S0(n369), .Y(n2127) );
  MXI2XL U759 ( .A(n888), .B(n3695), .S0(n369), .Y(n2128) );
  MXI2XL U760 ( .A(n889), .B(n3694), .S0(n369), .Y(n2129) );
  MXI2XL U761 ( .A(n890), .B(n3693), .S0(n370), .Y(n2130) );
  MXI2XL U762 ( .A(n891), .B(n3692), .S0(n370), .Y(n2131) );
  MXI2XL U763 ( .A(n892), .B(n3691), .S0(n370), .Y(n2132) );
  MXI2XL U764 ( .A(n893), .B(n3690), .S0(n370), .Y(n2133) );
  MXI2XL U765 ( .A(n894), .B(n3689), .S0(n370), .Y(n2134) );
  MXI2XL U766 ( .A(n895), .B(n3688), .S0(n370), .Y(n2135) );
  MXI2XL U767 ( .A(n896), .B(n3687), .S0(n370), .Y(n2136) );
  MXI2XL U768 ( .A(n897), .B(n3686), .S0(n370), .Y(n2137) );
  MXI2XL U769 ( .A(n898), .B(n3685), .S0(n370), .Y(n2138) );
  MXI2XL U770 ( .A(n899), .B(n3684), .S0(n370), .Y(n2139) );
  MXI2XL U771 ( .A(n900), .B(n3683), .S0(n370), .Y(n2140) );
  MXI2XL U772 ( .A(n901), .B(n3682), .S0(n370), .Y(n2141) );
  MXI2XL U773 ( .A(n902), .B(n3681), .S0(n370), .Y(n2142) );
  MXI2XL U774 ( .A(n903), .B(n3680), .S0(n371), .Y(n2143) );
  MXI2XL U775 ( .A(n904), .B(n3679), .S0(n371), .Y(n2144) );
  MXI2XL U776 ( .A(n905), .B(n3678), .S0(n371), .Y(n2145) );
  MXI2XL U777 ( .A(n906), .B(n3677), .S0(n371), .Y(n2146) );
  MXI2XL U778 ( .A(n907), .B(n3676), .S0(n371), .Y(n2147) );
  MXI2XL U779 ( .A(n908), .B(n3675), .S0(n371), .Y(n2148) );
  MXI2XL U780 ( .A(n909), .B(n3674), .S0(n371), .Y(n2149) );
  MXI2XL U781 ( .A(n910), .B(n3673), .S0(n371), .Y(n2150) );
  MXI2XL U782 ( .A(n911), .B(n3672), .S0(n371), .Y(n2151) );
  MXI2XL U783 ( .A(n912), .B(n3671), .S0(n371), .Y(n2152) );
  MXI2XL U784 ( .A(n913), .B(n3670), .S0(n371), .Y(n2153) );
  MXI2XL U785 ( .A(n914), .B(n3669), .S0(n371), .Y(n2154) );
  MXI2XL U786 ( .A(n947), .B(n3636), .S0(n3737), .Y(n2187) );
  MXI2XL U787 ( .A(n948), .B(n3635), .S0(n369), .Y(n2188) );
  MXI2XL U788 ( .A(n949), .B(n3634), .S0(n373), .Y(n2189) );
  MXI2XL U789 ( .A(n950), .B(n3633), .S0(n370), .Y(n2190) );
  MXI2XL U790 ( .A(n951), .B(n3632), .S0(n374), .Y(n2191) );
  MXI2XL U791 ( .A(n952), .B(n3631), .S0(n367), .Y(n2192) );
  MXI2XL U792 ( .A(n953), .B(n3630), .S0(n368), .Y(n2193) );
  MXI2XL U793 ( .A(n954), .B(n3629), .S0(n371), .Y(n2194) );
  MXI2XL U794 ( .A(n955), .B(n3628), .S0(n374), .Y(n2195) );
  MXI2XL U795 ( .A(n956), .B(n3627), .S0(n374), .Y(n2196) );
  MXI2XL U796 ( .A(n957), .B(n3626), .S0(n374), .Y(n2197) );
  MXI2XL U797 ( .A(n958), .B(n3625), .S0(n374), .Y(n2198) );
  MXI2XL U798 ( .A(n959), .B(n3624), .S0(n374), .Y(n2199) );
  MXI2XL U799 ( .A(n960), .B(n3623), .S0(n374), .Y(n2200) );
  MXI2XL U800 ( .A(n961), .B(n3622), .S0(n374), .Y(n2201) );
  MXI2XL U801 ( .A(n962), .B(n3621), .S0(n374), .Y(n2202) );
  MXI2XL U802 ( .A(n963), .B(n3620), .S0(n374), .Y(n2203) );
  MXI2XL U803 ( .A(n964), .B(n3619), .S0(n374), .Y(n2204) );
  MXI2XL U804 ( .A(n965), .B(n3618), .S0(n374), .Y(n2205) );
  MXI2XL U805 ( .A(n966), .B(n3617), .S0(n374), .Y(n2206) );
  MXI2XL U806 ( .A(n967), .B(n3616), .S0(n374), .Y(n2207) );
  MXI2XL U807 ( .A(n968), .B(n3615), .S0(n368), .Y(n2208) );
  MXI2XL U808 ( .A(n969), .B(n3614), .S0(n371), .Y(n2209) );
  MXI2XL U809 ( .A(n970), .B(n3613), .S0(n375), .Y(n2210) );
  MXI2XL U810 ( .A(n971), .B(n3612), .S0(n3737), .Y(n2211) );
  MXI2XL U811 ( .A(n972), .B(n3611), .S0(n372), .Y(n2212) );
  MXI2XL U812 ( .A(n973), .B(n3610), .S0(n369), .Y(n2213) );
  MXI2XL U813 ( .A(n974), .B(n3609), .S0(n373), .Y(n2214) );
  MXI2XL U814 ( .A(n975), .B(n3608), .S0(n370), .Y(n2215) );
  MXI2XL U815 ( .A(n976), .B(n3607), .S0(n374), .Y(n2216) );
  MXI2XL U816 ( .A(n977), .B(n3606), .S0(n367), .Y(n2217) );
  MXI2XL U817 ( .A(n978), .B(n3605), .S0(n368), .Y(n2218) );
  MXI2XL U818 ( .A(n1006), .B(n3732), .S0(n358), .Y(n2246) );
  MXI2XL U819 ( .A(n1007), .B(n3731), .S0(n358), .Y(n2247) );
  MXI2XL U820 ( .A(n1008), .B(n3730), .S0(n358), .Y(n2248) );
  MXI2XL U821 ( .A(n1009), .B(n3729), .S0(n358), .Y(n2249) );
  MXI2XL U822 ( .A(n1010), .B(n3728), .S0(n358), .Y(n2250) );
  MXI2XL U823 ( .A(n1011), .B(n3727), .S0(n358), .Y(n2251) );
  MXI2XL U824 ( .A(n1012), .B(n3726), .S0(n358), .Y(n2252) );
  MXI2XL U825 ( .A(n1013), .B(n3725), .S0(n358), .Y(n2253) );
  MXI2XL U826 ( .A(n1014), .B(n3724), .S0(n358), .Y(n2254) );
  MXI2XL U827 ( .A(n1015), .B(n3723), .S0(n358), .Y(n2255) );
  MXI2XL U828 ( .A(n1016), .B(n3722), .S0(n358), .Y(n2256) );
  MXI2XL U829 ( .A(n1017), .B(n3721), .S0(n358), .Y(n2257) );
  MXI2XL U830 ( .A(n1018), .B(n3720), .S0(n358), .Y(n2258) );
  MXI2XL U831 ( .A(n1019), .B(n3719), .S0(n359), .Y(n2259) );
  MXI2XL U832 ( .A(n1020), .B(n3718), .S0(n359), .Y(n2260) );
  MXI2XL U833 ( .A(n1021), .B(n3717), .S0(n359), .Y(n2261) );
  MXI2XL U834 ( .A(n1022), .B(n3716), .S0(n359), .Y(n2262) );
  MXI2XL U835 ( .A(n1023), .B(n3715), .S0(n359), .Y(n2263) );
  MXI2XL U836 ( .A(n1024), .B(n3714), .S0(n359), .Y(n2264) );
  MXI2XL U837 ( .A(n1025), .B(n3713), .S0(n359), .Y(n2265) );
  MXI2XL U838 ( .A(n1026), .B(n3712), .S0(n359), .Y(n2266) );
  MXI2XL U839 ( .A(n1027), .B(n3711), .S0(n359), .Y(n2267) );
  MXI2XL U840 ( .A(n1028), .B(n3710), .S0(n359), .Y(n2268) );
  MXI2XL U841 ( .A(n1029), .B(n3709), .S0(n359), .Y(n2269) );
  MXI2XL U842 ( .A(n1030), .B(n3708), .S0(n359), .Y(n2270) );
  MXI2XL U843 ( .A(n1031), .B(n3707), .S0(n359), .Y(n2271) );
  MXI2XL U844 ( .A(n1032), .B(n3706), .S0(n360), .Y(n2272) );
  MXI2XL U845 ( .A(n1033), .B(n3705), .S0(n360), .Y(n2273) );
  MXI2XL U846 ( .A(n1034), .B(n3704), .S0(n360), .Y(n2274) );
  MXI2XL U847 ( .A(n1035), .B(n3703), .S0(n360), .Y(n2275) );
  MXI2XL U848 ( .A(n1036), .B(n3702), .S0(n360), .Y(n2276) );
  MXI2XL U849 ( .A(n1037), .B(n3701), .S0(n360), .Y(n2277) );
  MXI2XL U850 ( .A(n1038), .B(n3700), .S0(n360), .Y(n2278) );
  MXI2XL U851 ( .A(n1039), .B(n3699), .S0(n360), .Y(n2279) );
  MXI2XL U852 ( .A(n1040), .B(n3698), .S0(n360), .Y(n2280) );
  MXI2XL U853 ( .A(n1041), .B(n3697), .S0(n360), .Y(n2281) );
  MXI2XL U854 ( .A(n1042), .B(n3696), .S0(n360), .Y(n2282) );
  MXI2XL U855 ( .A(n1043), .B(n3695), .S0(n360), .Y(n2283) );
  MXI2XL U856 ( .A(n1044), .B(n3694), .S0(n360), .Y(n2284) );
  MXI2XL U857 ( .A(n1045), .B(n3693), .S0(n361), .Y(n2285) );
  MXI2XL U858 ( .A(n1046), .B(n3692), .S0(n361), .Y(n2286) );
  MXI2XL U859 ( .A(n1047), .B(n3691), .S0(n361), .Y(n2287) );
  MXI2XL U860 ( .A(n1048), .B(n3690), .S0(n361), .Y(n2288) );
  MXI2XL U861 ( .A(n1049), .B(n3689), .S0(n361), .Y(n2289) );
  MXI2XL U862 ( .A(n1050), .B(n3688), .S0(n361), .Y(n2290) );
  MXI2XL U863 ( .A(n1051), .B(n3687), .S0(n361), .Y(n2291) );
  MXI2XL U864 ( .A(n1052), .B(n3686), .S0(n361), .Y(n2292) );
  MXI2XL U865 ( .A(n1053), .B(n3685), .S0(n361), .Y(n2293) );
  MXI2XL U866 ( .A(n1054), .B(n3684), .S0(n361), .Y(n2294) );
  MXI2XL U867 ( .A(n1055), .B(n3683), .S0(n361), .Y(n2295) );
  MXI2XL U868 ( .A(n1056), .B(n3682), .S0(n361), .Y(n2296) );
  MXI2XL U869 ( .A(n1057), .B(n3681), .S0(n361), .Y(n2297) );
  MXI2XL U870 ( .A(n1058), .B(n3680), .S0(n362), .Y(n2298) );
  MXI2XL U871 ( .A(n1059), .B(n3679), .S0(n362), .Y(n2299) );
  MXI2XL U872 ( .A(n1060), .B(n3678), .S0(n362), .Y(n2300) );
  MXI2XL U873 ( .A(n1061), .B(n3677), .S0(n362), .Y(n2301) );
  MXI2XL U874 ( .A(n1062), .B(n3676), .S0(n362), .Y(n2302) );
  MXI2XL U875 ( .A(n1063), .B(n3675), .S0(n362), .Y(n2303) );
  MXI2XL U876 ( .A(n1064), .B(n3674), .S0(n362), .Y(n2304) );
  MXI2XL U877 ( .A(n1065), .B(n3673), .S0(n362), .Y(n2305) );
  MXI2XL U878 ( .A(n1066), .B(n3672), .S0(n362), .Y(n2306) );
  MXI2XL U879 ( .A(n1067), .B(n3671), .S0(n362), .Y(n2307) );
  MXI2XL U880 ( .A(n1068), .B(n3670), .S0(n362), .Y(n2308) );
  MXI2XL U881 ( .A(n1069), .B(n3669), .S0(n362), .Y(n2309) );
  MXI2XL U882 ( .A(n1102), .B(n3636), .S0(n3736), .Y(n2342) );
  MXI2XL U883 ( .A(n1103), .B(n3635), .S0(n360), .Y(n2343) );
  MXI2XL U884 ( .A(n1104), .B(n3634), .S0(n364), .Y(n2344) );
  MXI2XL U885 ( .A(n1105), .B(n3633), .S0(n361), .Y(n2345) );
  MXI2XL U886 ( .A(n1106), .B(n3632), .S0(n365), .Y(n2346) );
  MXI2XL U887 ( .A(n1107), .B(n3631), .S0(n358), .Y(n2347) );
  MXI2XL U888 ( .A(n1108), .B(n3630), .S0(n359), .Y(n2348) );
  MXI2XL U889 ( .A(n1109), .B(n3629), .S0(n362), .Y(n2349) );
  MXI2XL U890 ( .A(n1110), .B(n3628), .S0(n365), .Y(n2350) );
  MXI2XL U891 ( .A(n1111), .B(n3627), .S0(n365), .Y(n2351) );
  MXI2XL U892 ( .A(n1112), .B(n3626), .S0(n365), .Y(n2352) );
  MXI2XL U893 ( .A(n1113), .B(n3625), .S0(n365), .Y(n2353) );
  MXI2XL U894 ( .A(n1114), .B(n3624), .S0(n365), .Y(n2354) );
  MXI2XL U895 ( .A(n1115), .B(n3623), .S0(n365), .Y(n2355) );
  MXI2XL U896 ( .A(n1116), .B(n3622), .S0(n365), .Y(n2356) );
  MXI2XL U897 ( .A(n1117), .B(n3621), .S0(n365), .Y(n2357) );
  MXI2XL U898 ( .A(n1118), .B(n3620), .S0(n365), .Y(n2358) );
  MXI2XL U899 ( .A(n1119), .B(n3619), .S0(n365), .Y(n2359) );
  MXI2XL U900 ( .A(n1120), .B(n3618), .S0(n365), .Y(n2360) );
  MXI2XL U901 ( .A(n1121), .B(n3617), .S0(n365), .Y(n2361) );
  MXI2XL U902 ( .A(n1122), .B(n3616), .S0(n365), .Y(n2362) );
  MXI2XL U903 ( .A(n1123), .B(n3615), .S0(n359), .Y(n2363) );
  MXI2XL U904 ( .A(n1124), .B(n3614), .S0(n362), .Y(n2364) );
  MXI2XL U905 ( .A(n1125), .B(n3613), .S0(n366), .Y(n2365) );
  MXI2XL U906 ( .A(n1126), .B(n3612), .S0(n3736), .Y(n2366) );
  MXI2XL U907 ( .A(n1127), .B(n3611), .S0(n363), .Y(n2367) );
  MXI2XL U908 ( .A(n1128), .B(n3610), .S0(n360), .Y(n2368) );
  MXI2XL U909 ( .A(n1129), .B(n3609), .S0(n364), .Y(n2369) );
  MXI2XL U910 ( .A(n1130), .B(n3608), .S0(n361), .Y(n2370) );
  MXI2XL U911 ( .A(n1131), .B(n3607), .S0(n365), .Y(n2371) );
  MXI2XL U912 ( .A(n1132), .B(n3606), .S0(n358), .Y(n2372) );
  MXI2XL U913 ( .A(n1133), .B(n3605), .S0(n359), .Y(n2373) );
  MXI2XL U914 ( .A(n1161), .B(n3732), .S0(n349), .Y(n2401) );
  MXI2XL U915 ( .A(n1162), .B(n3731), .S0(n349), .Y(n2402) );
  MXI2XL U916 ( .A(n1163), .B(n3730), .S0(n349), .Y(n2403) );
  MXI2XL U917 ( .A(n1164), .B(n3729), .S0(n349), .Y(n2404) );
  MXI2XL U918 ( .A(n1165), .B(n3728), .S0(n349), .Y(n2405) );
  MXI2XL U919 ( .A(n1166), .B(n3727), .S0(n349), .Y(n2406) );
  MXI2XL U920 ( .A(n1167), .B(n3726), .S0(n349), .Y(n2407) );
  MXI2XL U921 ( .A(n1168), .B(n3725), .S0(n349), .Y(n2408) );
  MXI2XL U922 ( .A(n1169), .B(n3724), .S0(n349), .Y(n2409) );
  MXI2XL U923 ( .A(n1170), .B(n3723), .S0(n349), .Y(n2410) );
  MXI2XL U924 ( .A(n1171), .B(n3722), .S0(n349), .Y(n2411) );
  MXI2XL U925 ( .A(n1172), .B(n3721), .S0(n349), .Y(n2412) );
  MXI2XL U926 ( .A(n1173), .B(n3720), .S0(n349), .Y(n2413) );
  MXI2XL U927 ( .A(n1174), .B(n3719), .S0(n350), .Y(n2414) );
  MXI2XL U928 ( .A(n1175), .B(n3718), .S0(n350), .Y(n2415) );
  MXI2XL U929 ( .A(n1176), .B(n3717), .S0(n350), .Y(n2416) );
  MXI2XL U930 ( .A(n1177), .B(n3716), .S0(n350), .Y(n2417) );
  MXI2XL U931 ( .A(n1178), .B(n3715), .S0(n350), .Y(n2418) );
  MXI2XL U932 ( .A(n1179), .B(n3714), .S0(n350), .Y(n2419) );
  MXI2XL U933 ( .A(n1180), .B(n3713), .S0(n350), .Y(n2420) );
  MXI2XL U934 ( .A(n1181), .B(n3712), .S0(n350), .Y(n2421) );
  MXI2XL U935 ( .A(n1182), .B(n3711), .S0(n350), .Y(n2422) );
  MXI2XL U936 ( .A(n1183), .B(n3710), .S0(n350), .Y(n2423) );
  MXI2XL U937 ( .A(n1184), .B(n3709), .S0(n350), .Y(n2424) );
  MXI2XL U938 ( .A(n1185), .B(n3708), .S0(n350), .Y(n2425) );
  MXI2XL U939 ( .A(n1186), .B(n3707), .S0(n350), .Y(n2426) );
  MXI2XL U940 ( .A(n1187), .B(n3706), .S0(n351), .Y(n2427) );
  MXI2XL U941 ( .A(n1188), .B(n3705), .S0(n351), .Y(n2428) );
  MXI2XL U942 ( .A(n1189), .B(n3704), .S0(n351), .Y(n2429) );
  MXI2XL U943 ( .A(n1190), .B(n3703), .S0(n351), .Y(n2430) );
  MXI2XL U944 ( .A(n1191), .B(n3702), .S0(n351), .Y(n2431) );
  MXI2XL U945 ( .A(n1192), .B(n3701), .S0(n351), .Y(n2432) );
  MXI2XL U946 ( .A(n1193), .B(n3700), .S0(n351), .Y(n2433) );
  MXI2XL U947 ( .A(n1194), .B(n3699), .S0(n351), .Y(n2434) );
  MXI2XL U948 ( .A(n1195), .B(n3698), .S0(n351), .Y(n2435) );
  MXI2XL U949 ( .A(n1196), .B(n3697), .S0(n351), .Y(n2436) );
  MXI2XL U950 ( .A(n1197), .B(n3696), .S0(n351), .Y(n2437) );
  MXI2XL U951 ( .A(n1198), .B(n3695), .S0(n351), .Y(n2438) );
  MXI2XL U952 ( .A(n1199), .B(n3694), .S0(n351), .Y(n2439) );
  MXI2XL U953 ( .A(n1200), .B(n3693), .S0(n352), .Y(n2440) );
  MXI2XL U954 ( .A(n1201), .B(n3692), .S0(n352), .Y(n2441) );
  MXI2XL U955 ( .A(n1202), .B(n3691), .S0(n352), .Y(n2442) );
  MXI2XL U956 ( .A(n1203), .B(n3690), .S0(n352), .Y(n2443) );
  MXI2XL U957 ( .A(n1204), .B(n3689), .S0(n352), .Y(n2444) );
  MXI2XL U958 ( .A(n1205), .B(n3688), .S0(n352), .Y(n2445) );
  MXI2XL U959 ( .A(n1206), .B(n3687), .S0(n352), .Y(n2446) );
  MXI2XL U960 ( .A(n1207), .B(n3686), .S0(n352), .Y(n2447) );
  MXI2XL U961 ( .A(n1208), .B(n3685), .S0(n352), .Y(n2448) );
  MXI2XL U962 ( .A(n1209), .B(n3684), .S0(n352), .Y(n2449) );
  MXI2XL U963 ( .A(n1210), .B(n3683), .S0(n352), .Y(n2450) );
  MXI2XL U964 ( .A(n1211), .B(n3682), .S0(n352), .Y(n2451) );
  MXI2XL U965 ( .A(n1212), .B(n3681), .S0(n352), .Y(n2452) );
  MXI2XL U966 ( .A(n1213), .B(n3680), .S0(n353), .Y(n2453) );
  MXI2XL U967 ( .A(n1214), .B(n3679), .S0(n353), .Y(n2454) );
  MXI2XL U968 ( .A(n1215), .B(n3678), .S0(n353), .Y(n2455) );
  MXI2XL U969 ( .A(n1216), .B(n3677), .S0(n353), .Y(n2456) );
  MXI2XL U970 ( .A(n1217), .B(n3676), .S0(n353), .Y(n2457) );
  MXI2XL U971 ( .A(n1218), .B(n3675), .S0(n353), .Y(n2458) );
  MXI2XL U972 ( .A(n1219), .B(n3674), .S0(n353), .Y(n2459) );
  MXI2XL U973 ( .A(n1220), .B(n3673), .S0(n353), .Y(n2460) );
  MXI2XL U974 ( .A(n1221), .B(n3672), .S0(n353), .Y(n2461) );
  MXI2XL U975 ( .A(n1222), .B(n3671), .S0(n353), .Y(n2462) );
  MXI2XL U976 ( .A(n1223), .B(n3670), .S0(n353), .Y(n2463) );
  MXI2XL U977 ( .A(n1224), .B(n3669), .S0(n353), .Y(n2464) );
  MXI2XL U978 ( .A(n1257), .B(n3636), .S0(n3735), .Y(n2497) );
  MXI2XL U979 ( .A(n1258), .B(n3635), .S0(n351), .Y(n2498) );
  MXI2XL U980 ( .A(n1259), .B(n3634), .S0(n355), .Y(n2499) );
  MXI2XL U981 ( .A(n1260), .B(n3633), .S0(n352), .Y(n2500) );
  MXI2XL U982 ( .A(n1261), .B(n3632), .S0(n356), .Y(n2501) );
  MXI2XL U983 ( .A(n1262), .B(n3631), .S0(n349), .Y(n2502) );
  MXI2XL U984 ( .A(n1263), .B(n3630), .S0(n350), .Y(n2503) );
  MXI2XL U985 ( .A(n1264), .B(n3629), .S0(n353), .Y(n2504) );
  MXI2XL U986 ( .A(n1265), .B(n3628), .S0(n356), .Y(n2505) );
  MXI2XL U987 ( .A(n1266), .B(n3627), .S0(n356), .Y(n2506) );
  MXI2XL U988 ( .A(n1267), .B(n3626), .S0(n356), .Y(n2507) );
  MXI2XL U989 ( .A(n1268), .B(n3625), .S0(n356), .Y(n2508) );
  MXI2XL U990 ( .A(n1269), .B(n3624), .S0(n356), .Y(n2509) );
  MXI2XL U991 ( .A(n1270), .B(n3623), .S0(n356), .Y(n2510) );
  MXI2XL U992 ( .A(n1271), .B(n3622), .S0(n356), .Y(n2511) );
  MXI2XL U993 ( .A(n1272), .B(n3621), .S0(n356), .Y(n2512) );
  MXI2XL U994 ( .A(n1273), .B(n3620), .S0(n356), .Y(n2513) );
  MXI2XL U995 ( .A(n1274), .B(n3619), .S0(n356), .Y(n2514) );
  MXI2XL U996 ( .A(n1275), .B(n3618), .S0(n356), .Y(n2515) );
  MXI2XL U997 ( .A(n1276), .B(n3617), .S0(n356), .Y(n2516) );
  MXI2XL U998 ( .A(n1277), .B(n3616), .S0(n356), .Y(n2517) );
  MXI2XL U999 ( .A(n1278), .B(n3615), .S0(n350), .Y(n2518) );
  MXI2XL U1000 ( .A(n1279), .B(n3614), .S0(n353), .Y(n2519) );
  MXI2XL U1001 ( .A(n1280), .B(n3613), .S0(n357), .Y(n2520) );
  MXI2XL U1002 ( .A(n1281), .B(n3612), .S0(n3735), .Y(n2521) );
  MXI2XL U1003 ( .A(n1282), .B(n3611), .S0(n354), .Y(n2522) );
  MXI2XL U1004 ( .A(n1283), .B(n3610), .S0(n351), .Y(n2523) );
  MXI2XL U1005 ( .A(n1284), .B(n3609), .S0(n355), .Y(n2524) );
  MXI2XL U1006 ( .A(n1285), .B(n3608), .S0(n352), .Y(n2525) );
  MXI2XL U1007 ( .A(n1286), .B(n3607), .S0(n356), .Y(n2526) );
  MXI2XL U1008 ( .A(n1287), .B(n3606), .S0(n349), .Y(n2527) );
  MXI2XL U1009 ( .A(n1288), .B(n3605), .S0(n350), .Y(n2528) );
  MXI2XL U1010 ( .A(n1316), .B(n3732), .S0(n340), .Y(n2556) );
  MXI2XL U1011 ( .A(n1317), .B(n3731), .S0(n340), .Y(n2557) );
  MXI2XL U1012 ( .A(n1318), .B(n3730), .S0(n340), .Y(n2558) );
  MXI2XL U1013 ( .A(n1319), .B(n3729), .S0(n340), .Y(n2559) );
  MXI2XL U1014 ( .A(n1320), .B(n3728), .S0(n340), .Y(n2560) );
  MXI2XL U1015 ( .A(n1321), .B(n3727), .S0(n340), .Y(n2561) );
  MXI2XL U1016 ( .A(n1322), .B(n3726), .S0(n340), .Y(n2562) );
  MXI2XL U1017 ( .A(n1323), .B(n3725), .S0(n340), .Y(n2563) );
  MXI2XL U1018 ( .A(n1324), .B(n3724), .S0(n340), .Y(n2564) );
  MXI2XL U1019 ( .A(n1325), .B(n3723), .S0(n340), .Y(n2565) );
  MXI2XL U1020 ( .A(n1326), .B(n3722), .S0(n340), .Y(n2566) );
  MXI2XL U1021 ( .A(n1327), .B(n3721), .S0(n340), .Y(n2567) );
  MXI2XL U1022 ( .A(n1328), .B(n3720), .S0(n340), .Y(n2568) );
  MXI2XL U1023 ( .A(n1329), .B(n3719), .S0(n341), .Y(n2569) );
  MXI2XL U1024 ( .A(n1330), .B(n3718), .S0(n341), .Y(n2570) );
  MXI2XL U1025 ( .A(n1331), .B(n3717), .S0(n341), .Y(n2571) );
  MXI2XL U1026 ( .A(n1332), .B(n3716), .S0(n341), .Y(n2572) );
  MXI2XL U1027 ( .A(n1333), .B(n3715), .S0(n341), .Y(n2573) );
  MXI2XL U1028 ( .A(n1334), .B(n3714), .S0(n341), .Y(n2574) );
  MXI2XL U1029 ( .A(n1335), .B(n3713), .S0(n341), .Y(n2575) );
  MXI2XL U1030 ( .A(n1336), .B(n3712), .S0(n341), .Y(n2576) );
  MXI2XL U1031 ( .A(n1337), .B(n3711), .S0(n341), .Y(n2577) );
  MXI2XL U1032 ( .A(n1338), .B(n3710), .S0(n341), .Y(n2578) );
  MXI2XL U1033 ( .A(n1339), .B(n3709), .S0(n341), .Y(n2579) );
  MXI2XL U1034 ( .A(n1340), .B(n3708), .S0(n341), .Y(n2580) );
  MXI2XL U1035 ( .A(n1341), .B(n3707), .S0(n341), .Y(n2581) );
  MXI2XL U1036 ( .A(n1342), .B(n3706), .S0(n342), .Y(n2582) );
  MXI2XL U1037 ( .A(n1343), .B(n3705), .S0(n342), .Y(n2583) );
  MXI2XL U1038 ( .A(n1344), .B(n3704), .S0(n342), .Y(n2584) );
  MXI2XL U1039 ( .A(n1345), .B(n3703), .S0(n342), .Y(n2585) );
  MXI2XL U1040 ( .A(n1346), .B(n3702), .S0(n342), .Y(n2586) );
  MXI2XL U1041 ( .A(n1347), .B(n3701), .S0(n342), .Y(n2587) );
  MXI2XL U1042 ( .A(n1348), .B(n3700), .S0(n342), .Y(n2588) );
  MXI2XL U1043 ( .A(n1349), .B(n3699), .S0(n342), .Y(n2589) );
  MXI2XL U1044 ( .A(n1350), .B(n3698), .S0(n342), .Y(n2590) );
  MXI2XL U1045 ( .A(n1351), .B(n3697), .S0(n342), .Y(n2591) );
  MXI2XL U1046 ( .A(n1352), .B(n3696), .S0(n342), .Y(n2592) );
  MXI2XL U1047 ( .A(n1353), .B(n3695), .S0(n342), .Y(n2593) );
  MXI2XL U1048 ( .A(n1354), .B(n3694), .S0(n342), .Y(n2594) );
  MXI2XL U1049 ( .A(n1355), .B(n3693), .S0(n343), .Y(n2595) );
  MXI2XL U1050 ( .A(n1356), .B(n3692), .S0(n343), .Y(n2596) );
  MXI2XL U1051 ( .A(n1357), .B(n3691), .S0(n343), .Y(n2597) );
  MXI2XL U1052 ( .A(n1358), .B(n3690), .S0(n343), .Y(n2598) );
  MXI2XL U1053 ( .A(n1359), .B(n3689), .S0(n343), .Y(n2599) );
  MXI2XL U1054 ( .A(n1360), .B(n3688), .S0(n343), .Y(n2600) );
  MXI2XL U1055 ( .A(n1361), .B(n3687), .S0(n343), .Y(n2601) );
  MXI2XL U1056 ( .A(n1362), .B(n3686), .S0(n343), .Y(n2602) );
  MXI2XL U1057 ( .A(n1363), .B(n3685), .S0(n343), .Y(n2603) );
  MXI2XL U1058 ( .A(n1364), .B(n3684), .S0(n343), .Y(n2604) );
  MXI2XL U1059 ( .A(n1365), .B(n3683), .S0(n343), .Y(n2605) );
  MXI2XL U1060 ( .A(n1366), .B(n3682), .S0(n343), .Y(n2606) );
  MXI2XL U1061 ( .A(n1367), .B(n3681), .S0(n343), .Y(n2607) );
  MXI2XL U1062 ( .A(n1368), .B(n3680), .S0(n344), .Y(n2608) );
  MXI2XL U1063 ( .A(n1369), .B(n3679), .S0(n344), .Y(n2609) );
  MXI2XL U1064 ( .A(n1370), .B(n3678), .S0(n344), .Y(n2610) );
  MXI2XL U1065 ( .A(n1371), .B(n3677), .S0(n344), .Y(n2611) );
  MXI2XL U1066 ( .A(n1372), .B(n3676), .S0(n344), .Y(n2612) );
  MXI2XL U1067 ( .A(n1373), .B(n3675), .S0(n344), .Y(n2613) );
  MXI2XL U1068 ( .A(n1374), .B(n3674), .S0(n344), .Y(n2614) );
  MXI2XL U1069 ( .A(n1375), .B(n3673), .S0(n344), .Y(n2615) );
  MXI2XL U1070 ( .A(n1376), .B(n3672), .S0(n344), .Y(n2616) );
  MXI2XL U1071 ( .A(n1377), .B(n3671), .S0(n344), .Y(n2617) );
  MXI2XL U1072 ( .A(n1378), .B(n3670), .S0(n344), .Y(n2618) );
  MXI2XL U1073 ( .A(n1379), .B(n3669), .S0(n344), .Y(n2619) );
  MXI2XL U1074 ( .A(n1412), .B(n3636), .S0(n3734), .Y(n2652) );
  MXI2XL U1075 ( .A(n1413), .B(n3635), .S0(n342), .Y(n2653) );
  MXI2XL U1076 ( .A(n1414), .B(n3634), .S0(n346), .Y(n2654) );
  MXI2XL U1077 ( .A(n1415), .B(n3633), .S0(n343), .Y(n2655) );
  MXI2XL U1078 ( .A(n1416), .B(n3632), .S0(n347), .Y(n2656) );
  MXI2XL U1079 ( .A(n1417), .B(n3631), .S0(n340), .Y(n2657) );
  MXI2XL U1080 ( .A(n1418), .B(n3630), .S0(n341), .Y(n2658) );
  MXI2XL U1081 ( .A(n1419), .B(n3629), .S0(n344), .Y(n2659) );
  MXI2XL U1082 ( .A(n1420), .B(n3628), .S0(n347), .Y(n2660) );
  MXI2XL U1083 ( .A(n1421), .B(n3627), .S0(n347), .Y(n2661) );
  MXI2XL U1084 ( .A(n1422), .B(n3626), .S0(n347), .Y(n2662) );
  MXI2XL U1085 ( .A(n1423), .B(n3625), .S0(n347), .Y(n2663) );
  MXI2XL U1086 ( .A(n1424), .B(n3624), .S0(n347), .Y(n2664) );
  MXI2XL U1087 ( .A(n1425), .B(n3623), .S0(n347), .Y(n2665) );
  MXI2XL U1088 ( .A(n1426), .B(n3622), .S0(n347), .Y(n2666) );
  MXI2XL U1089 ( .A(n1427), .B(n3621), .S0(n347), .Y(n2667) );
  MXI2XL U1090 ( .A(n1428), .B(n3620), .S0(n347), .Y(n2668) );
  MXI2XL U1091 ( .A(n1429), .B(n3619), .S0(n347), .Y(n2669) );
  MXI2XL U1092 ( .A(n1430), .B(n3618), .S0(n347), .Y(n2670) );
  MXI2XL U1093 ( .A(n1431), .B(n3617), .S0(n347), .Y(n2671) );
  MXI2XL U1094 ( .A(n1432), .B(n3616), .S0(n347), .Y(n2672) );
  MXI2XL U1095 ( .A(n1433), .B(n3615), .S0(n341), .Y(n2673) );
  MXI2XL U1096 ( .A(n1434), .B(n3614), .S0(n344), .Y(n2674) );
  MXI2XL U1097 ( .A(n1435), .B(n3613), .S0(n348), .Y(n2675) );
  MXI2XL U1098 ( .A(n1436), .B(n3612), .S0(n3734), .Y(n2676) );
  MXI2XL U1099 ( .A(n1437), .B(n3611), .S0(n345), .Y(n2677) );
  MXI2XL U1100 ( .A(n1438), .B(n3610), .S0(n342), .Y(n2678) );
  MXI2XL U1101 ( .A(n1439), .B(n3609), .S0(n346), .Y(n2679) );
  MXI2XL U1102 ( .A(n1440), .B(n3608), .S0(n343), .Y(n2680) );
  MXI2XL U1103 ( .A(n1441), .B(n3607), .S0(n347), .Y(n2681) );
  MXI2XL U1104 ( .A(n1442), .B(n3606), .S0(n340), .Y(n2682) );
  MXI2XL U1105 ( .A(n1443), .B(n3605), .S0(n341), .Y(n2683) );
  MXI2XL U1106 ( .A(n1471), .B(n3732), .S0(n331), .Y(n2711) );
  MXI2XL U1107 ( .A(n1472), .B(n3731), .S0(n331), .Y(n2712) );
  MXI2XL U1108 ( .A(n1473), .B(n3730), .S0(n331), .Y(n2713) );
  MXI2XL U1109 ( .A(n1474), .B(n3729), .S0(n331), .Y(n2714) );
  MXI2XL U1110 ( .A(n1475), .B(n3728), .S0(n331), .Y(n2715) );
  MXI2XL U1111 ( .A(n1476), .B(n3727), .S0(n331), .Y(n2716) );
  MXI2XL U1112 ( .A(n1477), .B(n3726), .S0(n331), .Y(n2717) );
  MXI2XL U1113 ( .A(n1478), .B(n3725), .S0(n331), .Y(n2718) );
  MXI2XL U1114 ( .A(n1479), .B(n3724), .S0(n331), .Y(n2719) );
  MXI2XL U1115 ( .A(n1480), .B(n3723), .S0(n331), .Y(n2720) );
  MXI2XL U1116 ( .A(n1481), .B(n3722), .S0(n331), .Y(n2721) );
  MXI2XL U1117 ( .A(n1482), .B(n3721), .S0(n331), .Y(n2722) );
  MXI2XL U1118 ( .A(n1483), .B(n3720), .S0(n331), .Y(n2723) );
  MXI2XL U1119 ( .A(n1484), .B(n3719), .S0(n332), .Y(n2724) );
  MXI2XL U1120 ( .A(n1485), .B(n3718), .S0(n332), .Y(n2725) );
  MXI2XL U1121 ( .A(n1486), .B(n3717), .S0(n332), .Y(n2726) );
  MXI2XL U1122 ( .A(n1487), .B(n3716), .S0(n332), .Y(n2727) );
  MXI2XL U1123 ( .A(n1488), .B(n3715), .S0(n332), .Y(n2728) );
  MXI2XL U1124 ( .A(n1489), .B(n3714), .S0(n332), .Y(n2729) );
  MXI2XL U1125 ( .A(n1490), .B(n3713), .S0(n332), .Y(n2730) );
  MXI2XL U1126 ( .A(n1491), .B(n3712), .S0(n332), .Y(n2731) );
  MXI2XL U1127 ( .A(n1492), .B(n3711), .S0(n332), .Y(n2732) );
  MXI2XL U1128 ( .A(n1493), .B(n3710), .S0(n332), .Y(n2733) );
  MXI2XL U1129 ( .A(n1494), .B(n3709), .S0(n332), .Y(n2734) );
  MXI2XL U1130 ( .A(n1495), .B(n3708), .S0(n332), .Y(n2735) );
  MXI2XL U1131 ( .A(n1496), .B(n3707), .S0(n332), .Y(n2736) );
  MXI2XL U1132 ( .A(n1497), .B(n3706), .S0(n333), .Y(n2737) );
  MXI2XL U1133 ( .A(n1498), .B(n3705), .S0(n333), .Y(n2738) );
  MXI2XL U1134 ( .A(n1499), .B(n3704), .S0(n333), .Y(n2739) );
  MXI2XL U1135 ( .A(n1500), .B(n3703), .S0(n333), .Y(n2740) );
  MXI2XL U1136 ( .A(n1501), .B(n3702), .S0(n333), .Y(n2741) );
  MXI2XL U1137 ( .A(n1502), .B(n3701), .S0(n333), .Y(n2742) );
  MXI2XL U1138 ( .A(n1503), .B(n3700), .S0(n333), .Y(n2743) );
  MXI2XL U1139 ( .A(n1504), .B(n3699), .S0(n333), .Y(n2744) );
  MXI2XL U1140 ( .A(n1505), .B(n3698), .S0(n333), .Y(n2745) );
  MXI2XL U1141 ( .A(n1506), .B(n3697), .S0(n333), .Y(n2746) );
  MXI2XL U1142 ( .A(n1507), .B(n3696), .S0(n333), .Y(n2747) );
  MXI2XL U1143 ( .A(n1508), .B(n3695), .S0(n333), .Y(n2748) );
  MXI2XL U1144 ( .A(n1509), .B(n3694), .S0(n333), .Y(n2749) );
  MXI2XL U1145 ( .A(n1510), .B(n3693), .S0(n334), .Y(n2750) );
  MXI2XL U1146 ( .A(n1511), .B(n3692), .S0(n334), .Y(n2751) );
  MXI2XL U1147 ( .A(n1512), .B(n3691), .S0(n334), .Y(n2752) );
  MXI2XL U1148 ( .A(n1513), .B(n3690), .S0(n334), .Y(n2753) );
  MXI2XL U1149 ( .A(n1514), .B(n3689), .S0(n334), .Y(n2754) );
  MXI2XL U1150 ( .A(n1515), .B(n3688), .S0(n334), .Y(n2755) );
  MXI2XL U1151 ( .A(n1516), .B(n3687), .S0(n334), .Y(n2756) );
  MXI2XL U1152 ( .A(n1517), .B(n3686), .S0(n334), .Y(n2757) );
  MXI2XL U1153 ( .A(n1518), .B(n3685), .S0(n334), .Y(n2758) );
  MXI2XL U1154 ( .A(n1519), .B(n3684), .S0(n334), .Y(n2759) );
  MXI2XL U1155 ( .A(n1520), .B(n3683), .S0(n334), .Y(n2760) );
  MXI2XL U1156 ( .A(n1521), .B(n3682), .S0(n334), .Y(n2761) );
  MXI2XL U1157 ( .A(n1522), .B(n3681), .S0(n334), .Y(n2762) );
  MXI2XL U1158 ( .A(n1523), .B(n3680), .S0(n335), .Y(n2763) );
  MXI2XL U1159 ( .A(n1524), .B(n3679), .S0(n335), .Y(n2764) );
  MXI2XL U1160 ( .A(n1525), .B(n3678), .S0(n335), .Y(n2765) );
  MXI2XL U1161 ( .A(n1526), .B(n3677), .S0(n335), .Y(n2766) );
  MXI2XL U1162 ( .A(n1527), .B(n3676), .S0(n335), .Y(n2767) );
  MXI2XL U1163 ( .A(n1528), .B(n3675), .S0(n335), .Y(n2768) );
  MXI2XL U1164 ( .A(n1529), .B(n3674), .S0(n335), .Y(n2769) );
  MXI2XL U1165 ( .A(n1530), .B(n3673), .S0(n335), .Y(n2770) );
  MXI2XL U1166 ( .A(n1531), .B(n3672), .S0(n335), .Y(n2771) );
  MXI2XL U1167 ( .A(n1532), .B(n3671), .S0(n335), .Y(n2772) );
  MXI2XL U1168 ( .A(n1533), .B(n3670), .S0(n335), .Y(n2773) );
  MXI2XL U1169 ( .A(n1534), .B(n3669), .S0(n335), .Y(n2774) );
  MXI2XL U1170 ( .A(n1567), .B(n3636), .S0(n3733), .Y(n2807) );
  MXI2XL U1171 ( .A(n1568), .B(n3635), .S0(n333), .Y(n2808) );
  MXI2XL U1172 ( .A(n1569), .B(n3634), .S0(n337), .Y(n2809) );
  MXI2XL U1173 ( .A(n1570), .B(n3633), .S0(n334), .Y(n2810) );
  MXI2XL U1174 ( .A(n1571), .B(n3632), .S0(n338), .Y(n2811) );
  MXI2XL U1175 ( .A(n1572), .B(n3631), .S0(n331), .Y(n2812) );
  MXI2XL U1176 ( .A(n1573), .B(n3630), .S0(n332), .Y(n2813) );
  MXI2XL U1177 ( .A(n1574), .B(n3629), .S0(n335), .Y(n2814) );
  MXI2XL U1178 ( .A(n1575), .B(n3628), .S0(n338), .Y(n2815) );
  MXI2XL U1179 ( .A(n1576), .B(n3627), .S0(n338), .Y(n2816) );
  MXI2XL U1180 ( .A(n1577), .B(n3626), .S0(n338), .Y(n2817) );
  MXI2XL U1181 ( .A(n1578), .B(n3625), .S0(n338), .Y(n2818) );
  MXI2XL U1182 ( .A(n1579), .B(n3624), .S0(n338), .Y(n2819) );
  MXI2XL U1183 ( .A(n1580), .B(n3623), .S0(n338), .Y(n2820) );
  MXI2XL U1184 ( .A(n1581), .B(n3622), .S0(n338), .Y(n2821) );
  MXI2XL U1185 ( .A(n1582), .B(n3621), .S0(n338), .Y(n2822) );
  MXI2XL U1186 ( .A(n1583), .B(n3620), .S0(n338), .Y(n2823) );
  MXI2XL U1187 ( .A(n1584), .B(n3619), .S0(n338), .Y(n2824) );
  MXI2XL U1188 ( .A(n1585), .B(n3618), .S0(n338), .Y(n2825) );
  MXI2XL U1189 ( .A(n1586), .B(n3617), .S0(n338), .Y(n2826) );
  MXI2XL U1190 ( .A(n1587), .B(n3616), .S0(n338), .Y(n2827) );
  MXI2XL U1191 ( .A(n1588), .B(n3615), .S0(n332), .Y(n2828) );
  MXI2XL U1192 ( .A(n1589), .B(n3614), .S0(n335), .Y(n2829) );
  MXI2XL U1193 ( .A(n1590), .B(n3613), .S0(n339), .Y(n2830) );
  MXI2XL U1194 ( .A(n1591), .B(n3612), .S0(n3733), .Y(n2831) );
  MXI2XL U1195 ( .A(n1592), .B(n3611), .S0(n336), .Y(n2832) );
  MXI2XL U1196 ( .A(n1593), .B(n3610), .S0(n333), .Y(n2833) );
  MXI2XL U1197 ( .A(n1594), .B(n3609), .S0(n337), .Y(n2834) );
  MXI2XL U1198 ( .A(n1595), .B(n3608), .S0(n334), .Y(n2835) );
  MXI2XL U1199 ( .A(n1596), .B(n3607), .S0(n338), .Y(n2836) );
  MXI2XL U1200 ( .A(n1597), .B(n3606), .S0(n331), .Y(n2837) );
  MXI2XL U1201 ( .A(n1598), .B(n3605), .S0(n332), .Y(n2838) );
  MXI2XL U1202 ( .A(n1626), .B(n3732), .S0(n322), .Y(n2866) );
  MXI2XL U1203 ( .A(n1627), .B(n3731), .S0(n322), .Y(n2867) );
  MXI2XL U1204 ( .A(n1628), .B(n3730), .S0(n322), .Y(n2868) );
  MXI2XL U1205 ( .A(n1629), .B(n3729), .S0(n322), .Y(n2869) );
  MXI2XL U1206 ( .A(n1630), .B(n3728), .S0(n322), .Y(n2870) );
  MXI2XL U1207 ( .A(n1631), .B(n3727), .S0(n322), .Y(n2871) );
  MXI2XL U1208 ( .A(n1632), .B(n3726), .S0(n322), .Y(n2872) );
  MXI2XL U1209 ( .A(n1633), .B(n3725), .S0(n322), .Y(n2873) );
  MXI2XL U1210 ( .A(n1634), .B(n3724), .S0(n322), .Y(n2874) );
  MXI2XL U1211 ( .A(n1635), .B(n3723), .S0(n322), .Y(n2875) );
  MXI2XL U1212 ( .A(n1636), .B(n3722), .S0(n322), .Y(n2876) );
  MXI2XL U1213 ( .A(n1637), .B(n3721), .S0(n322), .Y(n2877) );
  MXI2XL U1214 ( .A(n1638), .B(n3720), .S0(n322), .Y(n2878) );
  MXI2XL U1215 ( .A(n1639), .B(n3719), .S0(n323), .Y(n2879) );
  MXI2XL U1216 ( .A(n1640), .B(n3718), .S0(n323), .Y(n2880) );
  MXI2XL U1217 ( .A(n1641), .B(n3717), .S0(n323), .Y(n2881) );
  MXI2XL U1218 ( .A(n1642), .B(n3716), .S0(n323), .Y(n2882) );
  MXI2XL U1219 ( .A(n1643), .B(n3715), .S0(n323), .Y(n2883) );
  MXI2XL U1220 ( .A(n1644), .B(n3714), .S0(n323), .Y(n2884) );
  MXI2XL U1221 ( .A(n1645), .B(n3713), .S0(n323), .Y(n2885) );
  MXI2XL U1222 ( .A(n1646), .B(n3712), .S0(n323), .Y(n2886) );
  MXI2XL U1223 ( .A(n1647), .B(n3711), .S0(n323), .Y(n2887) );
  MXI2XL U1224 ( .A(n1648), .B(n3710), .S0(n323), .Y(n2888) );
  MXI2XL U1225 ( .A(n1649), .B(n3709), .S0(n323), .Y(n2889) );
  MXI2XL U1226 ( .A(n1650), .B(n3708), .S0(n323), .Y(n2890) );
  MXI2XL U1227 ( .A(n1651), .B(n3707), .S0(n323), .Y(n2891) );
  MXI2XL U1228 ( .A(n1652), .B(n3706), .S0(n324), .Y(n2892) );
  MXI2XL U1229 ( .A(n1653), .B(n3705), .S0(n324), .Y(n2893) );
  MXI2XL U1230 ( .A(n1654), .B(n3704), .S0(n324), .Y(n2894) );
  MXI2XL U1231 ( .A(n1655), .B(n3703), .S0(n324), .Y(n2895) );
  MXI2XL U1232 ( .A(n1656), .B(n3702), .S0(n324), .Y(n2896) );
  MXI2XL U1233 ( .A(n1657), .B(n3701), .S0(n324), .Y(n2897) );
  MXI2XL U1234 ( .A(n1658), .B(n3700), .S0(n324), .Y(n2898) );
  MXI2XL U1235 ( .A(n1659), .B(n3699), .S0(n324), .Y(n2899) );
  MXI2XL U1236 ( .A(n1660), .B(n3698), .S0(n324), .Y(n2900) );
  MXI2XL U1237 ( .A(n1661), .B(n3697), .S0(n324), .Y(n2901) );
  MXI2XL U1238 ( .A(n1662), .B(n3696), .S0(n324), .Y(n2902) );
  MXI2XL U1239 ( .A(n1663), .B(n3695), .S0(n324), .Y(n2903) );
  MXI2XL U1240 ( .A(n1664), .B(n3694), .S0(n324), .Y(n2904) );
  MXI2XL U1241 ( .A(n1665), .B(n3693), .S0(n325), .Y(n2905) );
  MXI2XL U1242 ( .A(n1666), .B(n3692), .S0(n325), .Y(n2906) );
  MXI2XL U1243 ( .A(n1667), .B(n3691), .S0(n325), .Y(n2907) );
  MXI2XL U1244 ( .A(n1668), .B(n3690), .S0(n325), .Y(n2908) );
  MXI2XL U1245 ( .A(n1669), .B(n3689), .S0(n325), .Y(n2909) );
  MXI2XL U1246 ( .A(n1670), .B(n3688), .S0(n325), .Y(n2910) );
  MXI2XL U1247 ( .A(n1671), .B(n3687), .S0(n325), .Y(n2911) );
  MXI2XL U1248 ( .A(n1672), .B(n3686), .S0(n325), .Y(n2912) );
  MXI2XL U1249 ( .A(n1673), .B(n3685), .S0(n325), .Y(n2913) );
  MXI2XL U1250 ( .A(n1674), .B(n3684), .S0(n325), .Y(n2914) );
  MXI2XL U1251 ( .A(n1675), .B(n3683), .S0(n325), .Y(n2915) );
  MXI2XL U1252 ( .A(n1676), .B(n3682), .S0(n325), .Y(n2916) );
  MXI2XL U1253 ( .A(n1677), .B(n3681), .S0(n325), .Y(n2917) );
  MXI2XL U1254 ( .A(n1678), .B(n3680), .S0(n326), .Y(n2918) );
  MXI2XL U1255 ( .A(n1679), .B(n3679), .S0(n326), .Y(n2919) );
  MXI2XL U1256 ( .A(n1680), .B(n3678), .S0(n326), .Y(n2920) );
  MXI2XL U1257 ( .A(n1681), .B(n3677), .S0(n326), .Y(n2921) );
  MXI2XL U1258 ( .A(n1682), .B(n3676), .S0(n326), .Y(n2922) );
  MXI2XL U1259 ( .A(n1683), .B(n3675), .S0(n326), .Y(n2923) );
  MXI2XL U1260 ( .A(n1684), .B(n3674), .S0(n326), .Y(n2924) );
  MXI2XL U1261 ( .A(n1685), .B(n3673), .S0(n326), .Y(n2925) );
  MXI2XL U1262 ( .A(n1686), .B(n3672), .S0(n326), .Y(n2926) );
  MXI2XL U1263 ( .A(n1687), .B(n3671), .S0(n326), .Y(n2927) );
  MXI2XL U1264 ( .A(n1688), .B(n3670), .S0(n326), .Y(n2928) );
  MXI2XL U1265 ( .A(n1689), .B(n3669), .S0(n326), .Y(n2929) );
  MXI2XL U1266 ( .A(n1722), .B(n3636), .S0(n3578), .Y(n2962) );
  MXI2XL U1267 ( .A(n1723), .B(n3635), .S0(n324), .Y(n2963) );
  MXI2XL U1268 ( .A(n1724), .B(n3634), .S0(n328), .Y(n2964) );
  MXI2XL U1269 ( .A(n1725), .B(n3633), .S0(n325), .Y(n2965) );
  MXI2XL U1270 ( .A(n1726), .B(n3632), .S0(n329), .Y(n2966) );
  MXI2XL U1271 ( .A(n1727), .B(n3631), .S0(n322), .Y(n2967) );
  MXI2XL U1272 ( .A(n1728), .B(n3630), .S0(n323), .Y(n2968) );
  MXI2XL U1273 ( .A(n1729), .B(n3629), .S0(n326), .Y(n2969) );
  MXI2XL U1274 ( .A(n1730), .B(n3628), .S0(n329), .Y(n2970) );
  MXI2XL U1275 ( .A(n1731), .B(n3627), .S0(n329), .Y(n2971) );
  MXI2XL U1276 ( .A(n1732), .B(n3626), .S0(n329), .Y(n2972) );
  MXI2XL U1277 ( .A(n1733), .B(n3625), .S0(n329), .Y(n2973) );
  MXI2XL U1278 ( .A(n1734), .B(n3624), .S0(n329), .Y(n2974) );
  MXI2XL U1279 ( .A(n1735), .B(n3623), .S0(n329), .Y(n2975) );
  MXI2XL U1280 ( .A(n1736), .B(n3622), .S0(n329), .Y(n2976) );
  MXI2XL U1281 ( .A(n1737), .B(n3621), .S0(n329), .Y(n2977) );
  MXI2XL U1282 ( .A(n1738), .B(n3620), .S0(n329), .Y(n2978) );
  MXI2XL U1283 ( .A(n1739), .B(n3619), .S0(n329), .Y(n2979) );
  MXI2XL U1284 ( .A(n1740), .B(n3618), .S0(n329), .Y(n2980) );
  MXI2XL U1285 ( .A(n1741), .B(n3617), .S0(n329), .Y(n2981) );
  MXI2XL U1286 ( .A(n1742), .B(n3616), .S0(n329), .Y(n2982) );
  MXI2XL U1287 ( .A(n1743), .B(n3615), .S0(n323), .Y(n2983) );
  MXI2XL U1288 ( .A(n1744), .B(n3614), .S0(n326), .Y(n2984) );
  MXI2XL U1289 ( .A(n1745), .B(n3613), .S0(n330), .Y(n2985) );
  MXI2XL U1290 ( .A(n1746), .B(n3612), .S0(n3578), .Y(n2986) );
  MXI2XL U1291 ( .A(n1747), .B(n3611), .S0(n327), .Y(n2987) );
  MXI2XL U1292 ( .A(n1748), .B(n3610), .S0(n324), .Y(n2988) );
  MXI2XL U1293 ( .A(n1749), .B(n3609), .S0(n328), .Y(n2989) );
  MXI2XL U1294 ( .A(n1750), .B(n3608), .S0(n325), .Y(n2990) );
  MXI2XL U1295 ( .A(n1751), .B(n3607), .S0(n329), .Y(n2991) );
  MXI2XL U1296 ( .A(n1752), .B(n3606), .S0(n322), .Y(n2992) );
  MXI2XL U1297 ( .A(n1753), .B(n3605), .S0(n323), .Y(n2993) );
  MXI2XL U1298 ( .A(n605), .B(n3668), .S0(n389), .Y(n1845) );
  MXI2XL U1299 ( .A(n606), .B(n3667), .S0(n390), .Y(n1846) );
  MXI2XL U1300 ( .A(n607), .B(n3666), .S0(n390), .Y(n1847) );
  MXI2XL U1301 ( .A(n608), .B(n3665), .S0(n390), .Y(n1848) );
  MXI2XL U1302 ( .A(n609), .B(n3664), .S0(n390), .Y(n1849) );
  MXI2XL U1303 ( .A(n610), .B(n3663), .S0(n390), .Y(n1850) );
  MXI2XL U1304 ( .A(n611), .B(n3662), .S0(n390), .Y(n1851) );
  MXI2XL U1305 ( .A(n612), .B(n3661), .S0(n390), .Y(n1852) );
  MXI2XL U1306 ( .A(n613), .B(n3660), .S0(n390), .Y(n1853) );
  MXI2XL U1307 ( .A(n614), .B(n3659), .S0(n390), .Y(n1854) );
  MXI2XL U1308 ( .A(n615), .B(n3658), .S0(n390), .Y(n1855) );
  MXI2XL U1309 ( .A(n616), .B(n3657), .S0(n390), .Y(n1856) );
  MXI2XL U1310 ( .A(n617), .B(n3656), .S0(n390), .Y(n1857) );
  MXI2XL U1311 ( .A(n618), .B(n3655), .S0(n390), .Y(n1858) );
  MXI2XL U1312 ( .A(n619), .B(n3654), .S0(n391), .Y(n1859) );
  MXI2XL U1313 ( .A(n620), .B(n3653), .S0(n391), .Y(n1860) );
  MXI2XL U1314 ( .A(n621), .B(n3652), .S0(n391), .Y(n1861) );
  MXI2XL U1315 ( .A(n622), .B(n3651), .S0(n391), .Y(n1862) );
  MXI2XL U1316 ( .A(n623), .B(n3650), .S0(n391), .Y(n1863) );
  MXI2XL U1317 ( .A(n624), .B(n3649), .S0(n391), .Y(n1864) );
  MXI2XL U1318 ( .A(n625), .B(n3648), .S0(n391), .Y(n1865) );
  MXI2XL U1319 ( .A(n626), .B(n3647), .S0(n391), .Y(n1866) );
  MXI2XL U1320 ( .A(n627), .B(n3646), .S0(n391), .Y(n1867) );
  MXI2XL U1321 ( .A(n628), .B(n3645), .S0(n391), .Y(n1868) );
  MXI2XL U1322 ( .A(n629), .B(n3644), .S0(n391), .Y(n1869) );
  MXI2XL U1323 ( .A(n630), .B(n3643), .S0(n391), .Y(n1870) );
  MXI2XL U1324 ( .A(n631), .B(n3642), .S0(n391), .Y(n1871) );
  MXI2XL U1325 ( .A(n632), .B(n3641), .S0(n385), .Y(n1872) );
  MXI2XL U1326 ( .A(n633), .B(n3640), .S0(n387), .Y(n1873) );
  MXI2XL U1327 ( .A(n634), .B(n3639), .S0(n391), .Y(n1874) );
  MXI2XL U1328 ( .A(n635), .B(n3638), .S0(n388), .Y(n1875) );
  MXI2XL U1329 ( .A(n636), .B(n3637), .S0(n392), .Y(n1876) );
  MXI2XL U1330 ( .A(n760), .B(n3668), .S0(n380), .Y(n2000) );
  MXI2XL U1331 ( .A(n761), .B(n3667), .S0(n381), .Y(n2001) );
  MXI2XL U1332 ( .A(n762), .B(n3666), .S0(n381), .Y(n2002) );
  MXI2XL U1333 ( .A(n763), .B(n3665), .S0(n381), .Y(n2003) );
  MXI2XL U1334 ( .A(n764), .B(n3664), .S0(n381), .Y(n2004) );
  MXI2XL U1335 ( .A(n765), .B(n3663), .S0(n381), .Y(n2005) );
  MXI2XL U1336 ( .A(n766), .B(n3662), .S0(n381), .Y(n2006) );
  MXI2XL U1337 ( .A(n767), .B(n3661), .S0(n381), .Y(n2007) );
  MXI2XL U1338 ( .A(n768), .B(n3660), .S0(n381), .Y(n2008) );
  MXI2XL U1339 ( .A(n769), .B(n3659), .S0(n381), .Y(n2009) );
  MXI2XL U1340 ( .A(n770), .B(n3658), .S0(n381), .Y(n2010) );
  MXI2XL U1341 ( .A(n771), .B(n3657), .S0(n381), .Y(n2011) );
  MXI2XL U1342 ( .A(n772), .B(n3656), .S0(n381), .Y(n2012) );
  MXI2XL U1343 ( .A(n773), .B(n3655), .S0(n381), .Y(n2013) );
  MXI2XL U1344 ( .A(n774), .B(n3654), .S0(n382), .Y(n2014) );
  MXI2XL U1345 ( .A(n775), .B(n3653), .S0(n382), .Y(n2015) );
  MXI2XL U1346 ( .A(n776), .B(n3652), .S0(n382), .Y(n2016) );
  MXI2XL U1347 ( .A(n777), .B(n3651), .S0(n382), .Y(n2017) );
  MXI2XL U1348 ( .A(n778), .B(n3650), .S0(n382), .Y(n2018) );
  MXI2XL U1349 ( .A(n779), .B(n3649), .S0(n382), .Y(n2019) );
  MXI2XL U1350 ( .A(n780), .B(n3648), .S0(n382), .Y(n2020) );
  MXI2XL U1351 ( .A(n781), .B(n3647), .S0(n382), .Y(n2021) );
  MXI2XL U1352 ( .A(n782), .B(n3646), .S0(n382), .Y(n2022) );
  MXI2XL U1353 ( .A(n783), .B(n3645), .S0(n382), .Y(n2023) );
  MXI2XL U1354 ( .A(n784), .B(n3644), .S0(n382), .Y(n2024) );
  MXI2XL U1355 ( .A(n785), .B(n3643), .S0(n382), .Y(n2025) );
  MXI2XL U1356 ( .A(n786), .B(n3642), .S0(n382), .Y(n2026) );
  MXI2XL U1357 ( .A(n787), .B(n3641), .S0(n376), .Y(n2027) );
  MXI2XL U1358 ( .A(n788), .B(n3640), .S0(n378), .Y(n2028) );
  MXI2XL U1359 ( .A(n789), .B(n3639), .S0(n382), .Y(n2029) );
  MXI2XL U1360 ( .A(n790), .B(n3638), .S0(n379), .Y(n2030) );
  MXI2XL U1361 ( .A(n791), .B(n3637), .S0(n383), .Y(n2031) );
  MXI2XL U1362 ( .A(n915), .B(n3668), .S0(n371), .Y(n2155) );
  MXI2XL U1363 ( .A(n916), .B(n3667), .S0(n372), .Y(n2156) );
  MXI2XL U1364 ( .A(n917), .B(n3666), .S0(n372), .Y(n2157) );
  MXI2XL U1365 ( .A(n918), .B(n3665), .S0(n372), .Y(n2158) );
  MXI2XL U1366 ( .A(n919), .B(n3664), .S0(n372), .Y(n2159) );
  MXI2XL U1367 ( .A(n920), .B(n3663), .S0(n372), .Y(n2160) );
  MXI2XL U1368 ( .A(n921), .B(n3662), .S0(n372), .Y(n2161) );
  MXI2XL U1369 ( .A(n922), .B(n3661), .S0(n372), .Y(n2162) );
  MXI2XL U1370 ( .A(n923), .B(n3660), .S0(n372), .Y(n2163) );
  MXI2XL U1371 ( .A(n924), .B(n3659), .S0(n372), .Y(n2164) );
  MXI2XL U1372 ( .A(n925), .B(n3658), .S0(n372), .Y(n2165) );
  MXI2XL U1373 ( .A(n926), .B(n3657), .S0(n372), .Y(n2166) );
  MXI2XL U1374 ( .A(n927), .B(n3656), .S0(n372), .Y(n2167) );
  MXI2XL U1375 ( .A(n928), .B(n3655), .S0(n372), .Y(n2168) );
  MXI2XL U1376 ( .A(n929), .B(n3654), .S0(n373), .Y(n2169) );
  MXI2XL U1377 ( .A(n930), .B(n3653), .S0(n373), .Y(n2170) );
  MXI2XL U1378 ( .A(n931), .B(n3652), .S0(n373), .Y(n2171) );
  MXI2XL U1379 ( .A(n932), .B(n3651), .S0(n373), .Y(n2172) );
  MXI2XL U1380 ( .A(n933), .B(n3650), .S0(n373), .Y(n2173) );
  MXI2XL U1381 ( .A(n934), .B(n3649), .S0(n373), .Y(n2174) );
  MXI2XL U1382 ( .A(n935), .B(n3648), .S0(n373), .Y(n2175) );
  MXI2XL U1383 ( .A(n936), .B(n3647), .S0(n373), .Y(n2176) );
  MXI2XL U1384 ( .A(n937), .B(n3646), .S0(n373), .Y(n2177) );
  MXI2XL U1385 ( .A(n938), .B(n3645), .S0(n373), .Y(n2178) );
  MXI2XL U1386 ( .A(n939), .B(n3644), .S0(n373), .Y(n2179) );
  MXI2XL U1387 ( .A(n940), .B(n3643), .S0(n373), .Y(n2180) );
  MXI2XL U1388 ( .A(n941), .B(n3642), .S0(n373), .Y(n2181) );
  MXI2XL U1389 ( .A(n942), .B(n3641), .S0(n367), .Y(n2182) );
  MXI2XL U1390 ( .A(n943), .B(n3640), .S0(n369), .Y(n2183) );
  MXI2XL U1391 ( .A(n944), .B(n3639), .S0(n373), .Y(n2184) );
  MXI2XL U1392 ( .A(n945), .B(n3638), .S0(n370), .Y(n2185) );
  MXI2XL U1393 ( .A(n946), .B(n3637), .S0(n374), .Y(n2186) );
  MXI2XL U1394 ( .A(n1070), .B(n3668), .S0(n362), .Y(n2310) );
  MXI2XL U1395 ( .A(n1071), .B(n3667), .S0(n363), .Y(n2311) );
  MXI2XL U1396 ( .A(n1072), .B(n3666), .S0(n363), .Y(n2312) );
  MXI2XL U1397 ( .A(n1073), .B(n3665), .S0(n363), .Y(n2313) );
  MXI2XL U1398 ( .A(n1074), .B(n3664), .S0(n363), .Y(n2314) );
  MXI2XL U1399 ( .A(n1075), .B(n3663), .S0(n363), .Y(n2315) );
  MXI2XL U1400 ( .A(n1076), .B(n3662), .S0(n363), .Y(n2316) );
  MXI2XL U1401 ( .A(n1077), .B(n3661), .S0(n363), .Y(n2317) );
  MXI2XL U1402 ( .A(n1078), .B(n3660), .S0(n363), .Y(n2318) );
  MXI2XL U1403 ( .A(n1079), .B(n3659), .S0(n363), .Y(n2319) );
  MXI2XL U1404 ( .A(n1080), .B(n3658), .S0(n363), .Y(n2320) );
  MXI2XL U1405 ( .A(n1081), .B(n3657), .S0(n363), .Y(n2321) );
  MXI2XL U1406 ( .A(n1082), .B(n3656), .S0(n363), .Y(n2322) );
  MXI2XL U1407 ( .A(n1083), .B(n3655), .S0(n363), .Y(n2323) );
  MXI2XL U1408 ( .A(n1084), .B(n3654), .S0(n364), .Y(n2324) );
  MXI2XL U1409 ( .A(n1085), .B(n3653), .S0(n364), .Y(n2325) );
  MXI2XL U1410 ( .A(n1086), .B(n3652), .S0(n364), .Y(n2326) );
  MXI2XL U1411 ( .A(n1087), .B(n3651), .S0(n364), .Y(n2327) );
  MXI2XL U1412 ( .A(n1088), .B(n3650), .S0(n364), .Y(n2328) );
  MXI2XL U1413 ( .A(n1089), .B(n3649), .S0(n364), .Y(n2329) );
  MXI2XL U1414 ( .A(n1090), .B(n3648), .S0(n364), .Y(n2330) );
  MXI2XL U1415 ( .A(n1091), .B(n3647), .S0(n364), .Y(n2331) );
  MXI2XL U1416 ( .A(n1092), .B(n3646), .S0(n364), .Y(n2332) );
  MXI2XL U1417 ( .A(n1093), .B(n3645), .S0(n364), .Y(n2333) );
  MXI2XL U1418 ( .A(n1094), .B(n3644), .S0(n364), .Y(n2334) );
  MXI2XL U1419 ( .A(n1095), .B(n3643), .S0(n364), .Y(n2335) );
  MXI2XL U1420 ( .A(n1096), .B(n3642), .S0(n364), .Y(n2336) );
  MXI2XL U1421 ( .A(n1097), .B(n3641), .S0(n358), .Y(n2337) );
  MXI2XL U1422 ( .A(n1098), .B(n3640), .S0(n360), .Y(n2338) );
  MXI2XL U1423 ( .A(n1099), .B(n3639), .S0(n364), .Y(n2339) );
  MXI2XL U1424 ( .A(n1100), .B(n3638), .S0(n361), .Y(n2340) );
  MXI2XL U1425 ( .A(n1101), .B(n3637), .S0(n365), .Y(n2341) );
  MXI2XL U1426 ( .A(n1225), .B(n3668), .S0(n353), .Y(n2465) );
  MXI2XL U1427 ( .A(n1226), .B(n3667), .S0(n354), .Y(n2466) );
  MXI2XL U1428 ( .A(n1227), .B(n3666), .S0(n354), .Y(n2467) );
  MXI2XL U1429 ( .A(n1228), .B(n3665), .S0(n354), .Y(n2468) );
  MXI2XL U1430 ( .A(n1229), .B(n3664), .S0(n354), .Y(n2469) );
  MXI2XL U1431 ( .A(n1230), .B(n3663), .S0(n354), .Y(n2470) );
  MXI2XL U1432 ( .A(n1231), .B(n3662), .S0(n354), .Y(n2471) );
  MXI2XL U1433 ( .A(n1232), .B(n3661), .S0(n354), .Y(n2472) );
  MXI2XL U1434 ( .A(n1233), .B(n3660), .S0(n354), .Y(n2473) );
  MXI2XL U1435 ( .A(n1234), .B(n3659), .S0(n354), .Y(n2474) );
  MXI2XL U1436 ( .A(n1235), .B(n3658), .S0(n354), .Y(n2475) );
  MXI2XL U1437 ( .A(n1236), .B(n3657), .S0(n354), .Y(n2476) );
  MXI2XL U1438 ( .A(n1237), .B(n3656), .S0(n354), .Y(n2477) );
  MXI2XL U1439 ( .A(n1238), .B(n3655), .S0(n354), .Y(n2478) );
  MXI2XL U1440 ( .A(n1239), .B(n3654), .S0(n355), .Y(n2479) );
  MXI2XL U1441 ( .A(n1240), .B(n3653), .S0(n355), .Y(n2480) );
  MXI2XL U1442 ( .A(n1241), .B(n3652), .S0(n355), .Y(n2481) );
  MXI2XL U1443 ( .A(n1242), .B(n3651), .S0(n355), .Y(n2482) );
  MXI2XL U1444 ( .A(n1243), .B(n3650), .S0(n355), .Y(n2483) );
  MXI2XL U1445 ( .A(n1244), .B(n3649), .S0(n355), .Y(n2484) );
  MXI2XL U1446 ( .A(n1245), .B(n3648), .S0(n355), .Y(n2485) );
  MXI2XL U1447 ( .A(n1246), .B(n3647), .S0(n355), .Y(n2486) );
  MXI2XL U1448 ( .A(n1247), .B(n3646), .S0(n355), .Y(n2487) );
  MXI2XL U1449 ( .A(n1248), .B(n3645), .S0(n355), .Y(n2488) );
  MXI2XL U1450 ( .A(n1249), .B(n3644), .S0(n355), .Y(n2489) );
  MXI2XL U1451 ( .A(n1250), .B(n3643), .S0(n355), .Y(n2490) );
  MXI2XL U1452 ( .A(n1251), .B(n3642), .S0(n355), .Y(n2491) );
  MXI2XL U1453 ( .A(n1252), .B(n3641), .S0(n349), .Y(n2492) );
  MXI2XL U1454 ( .A(n1253), .B(n3640), .S0(n351), .Y(n2493) );
  MXI2XL U1455 ( .A(n1254), .B(n3639), .S0(n355), .Y(n2494) );
  MXI2XL U1456 ( .A(n1255), .B(n3638), .S0(n352), .Y(n2495) );
  MXI2XL U1457 ( .A(n1256), .B(n3637), .S0(n356), .Y(n2496) );
  MXI2XL U1458 ( .A(n1380), .B(n3668), .S0(n344), .Y(n2620) );
  MXI2XL U1459 ( .A(n1381), .B(n3667), .S0(n345), .Y(n2621) );
  MXI2XL U1460 ( .A(n1382), .B(n3666), .S0(n345), .Y(n2622) );
  MXI2XL U1461 ( .A(n1383), .B(n3665), .S0(n345), .Y(n2623) );
  MXI2XL U1462 ( .A(n1384), .B(n3664), .S0(n345), .Y(n2624) );
  MXI2XL U1463 ( .A(n1385), .B(n3663), .S0(n345), .Y(n2625) );
  MXI2XL U1464 ( .A(n1386), .B(n3662), .S0(n345), .Y(n2626) );
  MXI2XL U1465 ( .A(n1387), .B(n3661), .S0(n345), .Y(n2627) );
  MXI2XL U1466 ( .A(n1388), .B(n3660), .S0(n345), .Y(n2628) );
  MXI2XL U1467 ( .A(n1389), .B(n3659), .S0(n345), .Y(n2629) );
  MXI2XL U1468 ( .A(n1390), .B(n3658), .S0(n345), .Y(n2630) );
  MXI2XL U1469 ( .A(n1391), .B(n3657), .S0(n345), .Y(n2631) );
  MXI2XL U1470 ( .A(n1392), .B(n3656), .S0(n345), .Y(n2632) );
  MXI2XL U1471 ( .A(n1393), .B(n3655), .S0(n345), .Y(n2633) );
  MXI2XL U1472 ( .A(n1394), .B(n3654), .S0(n346), .Y(n2634) );
  MXI2XL U1473 ( .A(n1395), .B(n3653), .S0(n346), .Y(n2635) );
  MXI2XL U1474 ( .A(n1396), .B(n3652), .S0(n346), .Y(n2636) );
  MXI2XL U1475 ( .A(n1397), .B(n3651), .S0(n346), .Y(n2637) );
  MXI2XL U1476 ( .A(n1398), .B(n3650), .S0(n346), .Y(n2638) );
  MXI2XL U1477 ( .A(n1399), .B(n3649), .S0(n346), .Y(n2639) );
  MXI2XL U1478 ( .A(n1400), .B(n3648), .S0(n346), .Y(n2640) );
  MXI2XL U1479 ( .A(n1401), .B(n3647), .S0(n346), .Y(n2641) );
  MXI2XL U1480 ( .A(n1402), .B(n3646), .S0(n346), .Y(n2642) );
  MXI2XL U1481 ( .A(n1403), .B(n3645), .S0(n346), .Y(n2643) );
  MXI2XL U1482 ( .A(n1404), .B(n3644), .S0(n346), .Y(n2644) );
  MXI2XL U1483 ( .A(n1405), .B(n3643), .S0(n346), .Y(n2645) );
  MXI2XL U1484 ( .A(n1406), .B(n3642), .S0(n346), .Y(n2646) );
  MXI2XL U1485 ( .A(n1407), .B(n3641), .S0(n340), .Y(n2647) );
  MXI2XL U1486 ( .A(n1408), .B(n3640), .S0(n342), .Y(n2648) );
  MXI2XL U1487 ( .A(n1409), .B(n3639), .S0(n346), .Y(n2649) );
  MXI2XL U1488 ( .A(n1410), .B(n3638), .S0(n343), .Y(n2650) );
  MXI2XL U1489 ( .A(n1411), .B(n3637), .S0(n347), .Y(n2651) );
  MXI2XL U1490 ( .A(n1535), .B(n3668), .S0(n335), .Y(n2775) );
  MXI2XL U1491 ( .A(n1536), .B(n3667), .S0(n336), .Y(n2776) );
  MXI2XL U1492 ( .A(n1537), .B(n3666), .S0(n336), .Y(n2777) );
  MXI2XL U1493 ( .A(n1538), .B(n3665), .S0(n336), .Y(n2778) );
  MXI2XL U1494 ( .A(n1539), .B(n3664), .S0(n336), .Y(n2779) );
  MXI2XL U1495 ( .A(n1540), .B(n3663), .S0(n336), .Y(n2780) );
  MXI2XL U1496 ( .A(n1541), .B(n3662), .S0(n336), .Y(n2781) );
  MXI2XL U1497 ( .A(n1542), .B(n3661), .S0(n336), .Y(n2782) );
  MXI2XL U1498 ( .A(n1543), .B(n3660), .S0(n336), .Y(n2783) );
  MXI2XL U1499 ( .A(n1544), .B(n3659), .S0(n336), .Y(n2784) );
  MXI2XL U1500 ( .A(n1545), .B(n3658), .S0(n336), .Y(n2785) );
  MXI2XL U1501 ( .A(n1546), .B(n3657), .S0(n336), .Y(n2786) );
  MXI2XL U1502 ( .A(n1547), .B(n3656), .S0(n336), .Y(n2787) );
  MXI2XL U1503 ( .A(n1548), .B(n3655), .S0(n336), .Y(n2788) );
  MXI2XL U1504 ( .A(n1549), .B(n3654), .S0(n337), .Y(n2789) );
  MXI2XL U1505 ( .A(n1550), .B(n3653), .S0(n337), .Y(n2790) );
  MXI2XL U1506 ( .A(n1551), .B(n3652), .S0(n337), .Y(n2791) );
  MXI2XL U1507 ( .A(n1552), .B(n3651), .S0(n337), .Y(n2792) );
  MXI2XL U1508 ( .A(n1553), .B(n3650), .S0(n337), .Y(n2793) );
  MXI2XL U1509 ( .A(n1554), .B(n3649), .S0(n337), .Y(n2794) );
  MXI2XL U1510 ( .A(n1555), .B(n3648), .S0(n337), .Y(n2795) );
  MXI2XL U1511 ( .A(n1556), .B(n3647), .S0(n337), .Y(n2796) );
  MXI2XL U1512 ( .A(n1557), .B(n3646), .S0(n337), .Y(n2797) );
  MXI2XL U1513 ( .A(n1558), .B(n3645), .S0(n337), .Y(n2798) );
  MXI2XL U1514 ( .A(n1559), .B(n3644), .S0(n337), .Y(n2799) );
  MXI2XL U1515 ( .A(n1560), .B(n3643), .S0(n337), .Y(n2800) );
  MXI2XL U1516 ( .A(n1561), .B(n3642), .S0(n337), .Y(n2801) );
  MXI2XL U1517 ( .A(n1562), .B(n3641), .S0(n331), .Y(n2802) );
  MXI2XL U1518 ( .A(n1563), .B(n3640), .S0(n333), .Y(n2803) );
  MXI2XL U1519 ( .A(n1564), .B(n3639), .S0(n337), .Y(n2804) );
  MXI2XL U1520 ( .A(n1565), .B(n3638), .S0(n334), .Y(n2805) );
  MXI2XL U1521 ( .A(n1566), .B(n3637), .S0(n338), .Y(n2806) );
  MXI2XL U1522 ( .A(n1690), .B(n3668), .S0(n326), .Y(n2930) );
  MXI2XL U1523 ( .A(n1691), .B(n3667), .S0(n327), .Y(n2931) );
  MXI2XL U1524 ( .A(n1692), .B(n3666), .S0(n327), .Y(n2932) );
  MXI2XL U1525 ( .A(n1693), .B(n3665), .S0(n327), .Y(n2933) );
  MXI2XL U1526 ( .A(n1694), .B(n3664), .S0(n327), .Y(n2934) );
  MXI2XL U1527 ( .A(n1695), .B(n3663), .S0(n327), .Y(n2935) );
  MXI2XL U1528 ( .A(n1696), .B(n3662), .S0(n327), .Y(n2936) );
  MXI2XL U1529 ( .A(n1697), .B(n3661), .S0(n327), .Y(n2937) );
  MXI2XL U1530 ( .A(n1698), .B(n3660), .S0(n327), .Y(n2938) );
  MXI2XL U1531 ( .A(n1699), .B(n3659), .S0(n327), .Y(n2939) );
  MXI2XL U1532 ( .A(n1700), .B(n3658), .S0(n327), .Y(n2940) );
  MXI2XL U1533 ( .A(n1701), .B(n3657), .S0(n327), .Y(n2941) );
  MXI2XL U1534 ( .A(n1702), .B(n3656), .S0(n327), .Y(n2942) );
  MXI2XL U1535 ( .A(n1703), .B(n3655), .S0(n327), .Y(n2943) );
  MXI2XL U1536 ( .A(n1704), .B(n3654), .S0(n328), .Y(n2944) );
  MXI2XL U1537 ( .A(n1705), .B(n3653), .S0(n328), .Y(n2945) );
  MXI2XL U1538 ( .A(n1706), .B(n3652), .S0(n328), .Y(n2946) );
  MXI2XL U1539 ( .A(n1707), .B(n3651), .S0(n328), .Y(n2947) );
  MXI2XL U1540 ( .A(n1708), .B(n3650), .S0(n328), .Y(n2948) );
  MXI2XL U1541 ( .A(n1709), .B(n3649), .S0(n328), .Y(n2949) );
  MXI2XL U1542 ( .A(n1710), .B(n3648), .S0(n328), .Y(n2950) );
  MXI2XL U1543 ( .A(n1711), .B(n3647), .S0(n328), .Y(n2951) );
  MXI2XL U1544 ( .A(n1712), .B(n3646), .S0(n328), .Y(n2952) );
  MXI2XL U1545 ( .A(n1713), .B(n3645), .S0(n328), .Y(n2953) );
  MXI2XL U1546 ( .A(n1714), .B(n3644), .S0(n328), .Y(n2954) );
  MXI2XL U1547 ( .A(n1715), .B(n3643), .S0(n328), .Y(n2955) );
  MXI2XL U1548 ( .A(n1716), .B(n3642), .S0(n328), .Y(n2956) );
  MXI2XL U1549 ( .A(n1717), .B(n3641), .S0(n322), .Y(n2957) );
  MXI2XL U1550 ( .A(n1718), .B(n3640), .S0(n324), .Y(n2958) );
  MXI2XL U1551 ( .A(n1719), .B(n3639), .S0(n328), .Y(n2959) );
  MXI2XL U1552 ( .A(n1720), .B(n3638), .S0(n325), .Y(n2960) );
  MXI2XL U1553 ( .A(n1721), .B(n3637), .S0(n329), .Y(n2961) );
  NAND2XL U1554 ( .A(proc_write), .B(n3764), .Y(n3762) );
  XOR2XL U1555 ( .A(proc_addr[17]), .B(N47), .Y(n3785) );
  XOR2XL U1556 ( .A(proc_addr[11]), .B(N53), .Y(n3792) );
  XOR2XL U1557 ( .A(proc_addr[23]), .B(N41), .Y(n3777) );
  XOR2XL U1558 ( .A(proc_addr[5]), .B(N59), .Y(n3799) );
  XOR2XL U1559 ( .A(proc_addr[18]), .B(N46), .Y(n3784) );
  XOR2XL U1560 ( .A(proc_addr[12]), .B(N52), .Y(n3791) );
  XOR2XL U1561 ( .A(proc_addr[24]), .B(N40), .Y(n3776) );
  XOR2XL U1562 ( .A(proc_addr[19]), .B(N45), .Y(n3786) );
  XOR2XL U1563 ( .A(proc_addr[13]), .B(N51), .Y(n3793) );
  XOR2XL U1564 ( .A(proc_addr[25]), .B(N39), .Y(n3778) );
  MXI2XL U1565 ( .A(n669), .B(n3604), .S0(n389), .Y(n1909) );
  MXI2XL U1566 ( .A(n670), .B(n3603), .S0(n393), .Y(n1910) );
  MXI2XL U1567 ( .A(n671), .B(n3602), .S0(n390), .Y(n1911) );
  MXI2XL U1568 ( .A(n672), .B(n3601), .S0(n388), .Y(n1912) );
  MXI2XL U1569 ( .A(n673), .B(n3600), .S0(n392), .Y(n1913) );
  MXI2XL U1570 ( .A(n674), .B(n3599), .S0(n385), .Y(n1914) );
  MXI2XL U1571 ( .A(n675), .B(n3598), .S0(n386), .Y(n1915) );
  MXI2XL U1572 ( .A(n676), .B(n3597), .S0(n389), .Y(n1916) );
  MXI2XL U1573 ( .A(n677), .B(n3596), .S0(n393), .Y(n1917) );
  MXI2XL U1574 ( .A(n678), .B(n3595), .S0(n390), .Y(n1918) );
  MXI2XL U1575 ( .A(n679), .B(n3594), .S0(n388), .Y(n1919) );
  MXI2XL U1576 ( .A(n680), .B(n3593), .S0(n392), .Y(n1920) );
  MXI2XL U1577 ( .A(n681), .B(n3592), .S0(n385), .Y(n1921) );
  MXI2XL U1578 ( .A(n682), .B(n3591), .S0(n386), .Y(n1922) );
  MXI2XL U1579 ( .A(n683), .B(n3590), .S0(n389), .Y(n1923) );
  MXI2XL U1580 ( .A(n684), .B(n3589), .S0(n393), .Y(n1924) );
  MXI2XL U1581 ( .A(n685), .B(n3588), .S0(n393), .Y(n1925) );
  MXI2XL U1582 ( .A(n686), .B(n3587), .S0(n393), .Y(n1926) );
  MXI2XL U1583 ( .A(n687), .B(n3586), .S0(n393), .Y(n1927) );
  MXI2XL U1584 ( .A(n688), .B(n3585), .S0(n393), .Y(n1928) );
  MXI2XL U1585 ( .A(n689), .B(n3584), .S0(n393), .Y(n1929) );
  MXI2XL U1586 ( .A(n690), .B(n3583), .S0(n393), .Y(n1930) );
  MXI2XL U1587 ( .A(n691), .B(n3582), .S0(n393), .Y(n1931) );
  MXI2XL U1588 ( .A(n692), .B(n3581), .S0(n393), .Y(n1932) );
  MXI2XL U1589 ( .A(n693), .B(n3580), .S0(n393), .Y(n1933) );
  MXI2XL U1590 ( .A(n824), .B(n3604), .S0(n380), .Y(n2064) );
  MXI2XL U1591 ( .A(n825), .B(n3603), .S0(n384), .Y(n2065) );
  MXI2XL U1592 ( .A(n826), .B(n3602), .S0(n381), .Y(n2066) );
  MXI2XL U1593 ( .A(n827), .B(n3601), .S0(n379), .Y(n2067) );
  MXI2XL U1594 ( .A(n828), .B(n3600), .S0(n383), .Y(n2068) );
  MXI2XL U1595 ( .A(n829), .B(n3599), .S0(n376), .Y(n2069) );
  MXI2XL U1596 ( .A(n830), .B(n3598), .S0(n377), .Y(n2070) );
  MXI2XL U1597 ( .A(n831), .B(n3597), .S0(n380), .Y(n2071) );
  MXI2XL U1598 ( .A(n832), .B(n3596), .S0(n384), .Y(n2072) );
  MXI2XL U1599 ( .A(n833), .B(n3595), .S0(n381), .Y(n2073) );
  MXI2XL U1600 ( .A(n834), .B(n3594), .S0(n379), .Y(n2074) );
  MXI2XL U1601 ( .A(n835), .B(n3593), .S0(n383), .Y(n2075) );
  MXI2XL U1602 ( .A(n836), .B(n3592), .S0(n376), .Y(n2076) );
  MXI2XL U1603 ( .A(n837), .B(n3591), .S0(n377), .Y(n2077) );
  MXI2XL U1604 ( .A(n838), .B(n3590), .S0(n380), .Y(n2078) );
  MXI2XL U1605 ( .A(n839), .B(n3589), .S0(n384), .Y(n2079) );
  MXI2XL U1606 ( .A(n840), .B(n3588), .S0(n384), .Y(n2080) );
  MXI2XL U1607 ( .A(n841), .B(n3587), .S0(n384), .Y(n2081) );
  MXI2XL U1608 ( .A(n842), .B(n3586), .S0(n384), .Y(n2082) );
  MXI2XL U1609 ( .A(n843), .B(n3585), .S0(n384), .Y(n2083) );
  MXI2XL U1610 ( .A(n844), .B(n3584), .S0(n384), .Y(n2084) );
  MXI2XL U1611 ( .A(n845), .B(n3583), .S0(n384), .Y(n2085) );
  MXI2XL U1612 ( .A(n846), .B(n3582), .S0(n384), .Y(n2086) );
  MXI2XL U1613 ( .A(n847), .B(n3581), .S0(n384), .Y(n2087) );
  MXI2XL U1614 ( .A(n848), .B(n3580), .S0(n384), .Y(n2088) );
  MXI2XL U1615 ( .A(n979), .B(n3604), .S0(n371), .Y(n2219) );
  MXI2XL U1616 ( .A(n980), .B(n3603), .S0(n375), .Y(n2220) );
  MXI2XL U1617 ( .A(n981), .B(n3602), .S0(n372), .Y(n2221) );
  MXI2XL U1618 ( .A(n982), .B(n3601), .S0(n370), .Y(n2222) );
  MXI2XL U1619 ( .A(n983), .B(n3600), .S0(n374), .Y(n2223) );
  MXI2XL U1620 ( .A(n984), .B(n3599), .S0(n367), .Y(n2224) );
  MXI2XL U1621 ( .A(n985), .B(n3598), .S0(n368), .Y(n2225) );
  MXI2XL U1622 ( .A(n986), .B(n3597), .S0(n371), .Y(n2226) );
  MXI2XL U1623 ( .A(n987), .B(n3596), .S0(n375), .Y(n2227) );
  MXI2XL U1624 ( .A(n988), .B(n3595), .S0(n372), .Y(n2228) );
  MXI2XL U1625 ( .A(n989), .B(n3594), .S0(n370), .Y(n2229) );
  MXI2XL U1626 ( .A(n990), .B(n3593), .S0(n374), .Y(n2230) );
  MXI2XL U1627 ( .A(n991), .B(n3592), .S0(n367), .Y(n2231) );
  MXI2XL U1628 ( .A(n992), .B(n3591), .S0(n368), .Y(n2232) );
  MXI2XL U1629 ( .A(n993), .B(n3590), .S0(n371), .Y(n2233) );
  MXI2XL U1630 ( .A(n994), .B(n3589), .S0(n375), .Y(n2234) );
  MXI2XL U1631 ( .A(n995), .B(n3588), .S0(n375), .Y(n2235) );
  MXI2XL U1632 ( .A(n996), .B(n3587), .S0(n375), .Y(n2236) );
  MXI2XL U1633 ( .A(n997), .B(n3586), .S0(n375), .Y(n2237) );
  MXI2XL U1634 ( .A(n998), .B(n3585), .S0(n375), .Y(n2238) );
  MXI2XL U1635 ( .A(n999), .B(n3584), .S0(n375), .Y(n2239) );
  MXI2XL U1636 ( .A(n1000), .B(n3583), .S0(n375), .Y(n2240) );
  MXI2XL U1637 ( .A(n1001), .B(n3582), .S0(n375), .Y(n2241) );
  MXI2XL U1638 ( .A(n1002), .B(n3581), .S0(n375), .Y(n2242) );
  MXI2XL U1639 ( .A(n1003), .B(n3580), .S0(n375), .Y(n2243) );
  MXI2XL U1640 ( .A(n1134), .B(n3604), .S0(n362), .Y(n2374) );
  MXI2XL U1641 ( .A(n1135), .B(n3603), .S0(n366), .Y(n2375) );
  MXI2XL U1642 ( .A(n1136), .B(n3602), .S0(n363), .Y(n2376) );
  MXI2XL U1643 ( .A(n1137), .B(n3601), .S0(n361), .Y(n2377) );
  MXI2XL U1644 ( .A(n1138), .B(n3600), .S0(n365), .Y(n2378) );
  MXI2XL U1645 ( .A(n1139), .B(n3599), .S0(n358), .Y(n2379) );
  MXI2XL U1646 ( .A(n1140), .B(n3598), .S0(n359), .Y(n2380) );
  MXI2XL U1647 ( .A(n1141), .B(n3597), .S0(n362), .Y(n2381) );
  MXI2XL U1648 ( .A(n1142), .B(n3596), .S0(n366), .Y(n2382) );
  MXI2XL U1649 ( .A(n1143), .B(n3595), .S0(n363), .Y(n2383) );
  MXI2XL U1650 ( .A(n1144), .B(n3594), .S0(n361), .Y(n2384) );
  MXI2XL U1651 ( .A(n1145), .B(n3593), .S0(n365), .Y(n2385) );
  MXI2XL U1652 ( .A(n1146), .B(n3592), .S0(n358), .Y(n2386) );
  MXI2XL U1653 ( .A(n1147), .B(n3591), .S0(n359), .Y(n2387) );
  MXI2XL U1654 ( .A(n1148), .B(n3590), .S0(n362), .Y(n2388) );
  MXI2XL U1655 ( .A(n1149), .B(n3589), .S0(n366), .Y(n2389) );
  MXI2XL U1656 ( .A(n1150), .B(n3588), .S0(n366), .Y(n2390) );
  MXI2XL U1657 ( .A(n1151), .B(n3587), .S0(n366), .Y(n2391) );
  MXI2XL U1658 ( .A(n1152), .B(n3586), .S0(n366), .Y(n2392) );
  MXI2XL U1659 ( .A(n1153), .B(n3585), .S0(n366), .Y(n2393) );
  MXI2XL U1660 ( .A(n1154), .B(n3584), .S0(n366), .Y(n2394) );
  MXI2XL U1661 ( .A(n1155), .B(n3583), .S0(n366), .Y(n2395) );
  MXI2XL U1662 ( .A(n1156), .B(n3582), .S0(n366), .Y(n2396) );
  MXI2XL U1663 ( .A(n1157), .B(n3581), .S0(n366), .Y(n2397) );
  MXI2XL U1664 ( .A(n1158), .B(n3580), .S0(n366), .Y(n2398) );
  MXI2XL U1665 ( .A(n1289), .B(n3604), .S0(n353), .Y(n2529) );
  MXI2XL U1666 ( .A(n1290), .B(n3603), .S0(n357), .Y(n2530) );
  MXI2XL U1667 ( .A(n1291), .B(n3602), .S0(n354), .Y(n2531) );
  MXI2XL U1668 ( .A(n1292), .B(n3601), .S0(n352), .Y(n2532) );
  MXI2XL U1669 ( .A(n1293), .B(n3600), .S0(n356), .Y(n2533) );
  MXI2XL U1670 ( .A(n1294), .B(n3599), .S0(n349), .Y(n2534) );
  MXI2XL U1671 ( .A(n1295), .B(n3598), .S0(n350), .Y(n2535) );
  MXI2XL U1672 ( .A(n1296), .B(n3597), .S0(n353), .Y(n2536) );
  MXI2XL U1673 ( .A(n1297), .B(n3596), .S0(n357), .Y(n2537) );
  MXI2XL U1674 ( .A(n1298), .B(n3595), .S0(n354), .Y(n2538) );
  MXI2XL U1675 ( .A(n1299), .B(n3594), .S0(n352), .Y(n2539) );
  MXI2XL U1676 ( .A(n1300), .B(n3593), .S0(n356), .Y(n2540) );
  MXI2XL U1677 ( .A(n1301), .B(n3592), .S0(n349), .Y(n2541) );
  MXI2XL U1678 ( .A(n1302), .B(n3591), .S0(n350), .Y(n2542) );
  MXI2XL U1679 ( .A(n1303), .B(n3590), .S0(n353), .Y(n2543) );
  MXI2XL U1680 ( .A(n1304), .B(n3589), .S0(n357), .Y(n2544) );
  MXI2XL U1681 ( .A(n1305), .B(n3588), .S0(n357), .Y(n2545) );
  MXI2XL U1682 ( .A(n1306), .B(n3587), .S0(n357), .Y(n2546) );
  MXI2XL U1683 ( .A(n1307), .B(n3586), .S0(n357), .Y(n2547) );
  MXI2XL U1684 ( .A(n1308), .B(n3585), .S0(n357), .Y(n2548) );
  MXI2XL U1685 ( .A(n1309), .B(n3584), .S0(n357), .Y(n2549) );
  MXI2XL U1686 ( .A(n1310), .B(n3583), .S0(n357), .Y(n2550) );
  MXI2XL U1687 ( .A(n1311), .B(n3582), .S0(n357), .Y(n2551) );
  MXI2XL U1688 ( .A(n1312), .B(n3581), .S0(n357), .Y(n2552) );
  MXI2XL U1689 ( .A(n1313), .B(n3580), .S0(n357), .Y(n2553) );
  MXI2XL U1690 ( .A(n1444), .B(n3604), .S0(n344), .Y(n2684) );
  MXI2XL U1691 ( .A(n1445), .B(n3603), .S0(n348), .Y(n2685) );
  MXI2XL U1692 ( .A(n1446), .B(n3602), .S0(n345), .Y(n2686) );
  MXI2XL U1693 ( .A(n1447), .B(n3601), .S0(n343), .Y(n2687) );
  MXI2XL U1694 ( .A(n1448), .B(n3600), .S0(n347), .Y(n2688) );
  MXI2XL U1695 ( .A(n1449), .B(n3599), .S0(n340), .Y(n2689) );
  MXI2XL U1696 ( .A(n1450), .B(n3598), .S0(n341), .Y(n2690) );
  MXI2XL U1697 ( .A(n1451), .B(n3597), .S0(n344), .Y(n2691) );
  MXI2XL U1698 ( .A(n1452), .B(n3596), .S0(n348), .Y(n2692) );
  MXI2XL U1699 ( .A(n1453), .B(n3595), .S0(n345), .Y(n2693) );
  MXI2XL U1700 ( .A(n1454), .B(n3594), .S0(n343), .Y(n2694) );
  MXI2XL U1701 ( .A(n1455), .B(n3593), .S0(n347), .Y(n2695) );
  MXI2XL U1702 ( .A(n1456), .B(n3592), .S0(n340), .Y(n2696) );
  MXI2XL U1703 ( .A(n1457), .B(n3591), .S0(n341), .Y(n2697) );
  MXI2XL U1704 ( .A(n1458), .B(n3590), .S0(n344), .Y(n2698) );
  MXI2XL U1705 ( .A(n1459), .B(n3589), .S0(n348), .Y(n2699) );
  MXI2XL U1706 ( .A(n1460), .B(n3588), .S0(n348), .Y(n2700) );
  MXI2XL U1707 ( .A(n1461), .B(n3587), .S0(n348), .Y(n2701) );
  MXI2XL U1708 ( .A(n1462), .B(n3586), .S0(n348), .Y(n2702) );
  MXI2XL U1709 ( .A(n1463), .B(n3585), .S0(n348), .Y(n2703) );
  MXI2XL U1710 ( .A(n1464), .B(n3584), .S0(n348), .Y(n2704) );
  MXI2XL U1711 ( .A(n1465), .B(n3583), .S0(n348), .Y(n2705) );
  MXI2XL U1712 ( .A(n1466), .B(n3582), .S0(n348), .Y(n2706) );
  MXI2XL U1713 ( .A(n1467), .B(n3581), .S0(n348), .Y(n2707) );
  MXI2XL U1714 ( .A(n1468), .B(n3580), .S0(n348), .Y(n2708) );
  MXI2XL U1715 ( .A(n1599), .B(n3604), .S0(n335), .Y(n2839) );
  MXI2XL U1716 ( .A(n1600), .B(n3603), .S0(n339), .Y(n2840) );
  MXI2XL U1717 ( .A(n1601), .B(n3602), .S0(n336), .Y(n2841) );
  MXI2XL U1718 ( .A(n1602), .B(n3601), .S0(n334), .Y(n2842) );
  MXI2XL U1719 ( .A(n1603), .B(n3600), .S0(n338), .Y(n2843) );
  MXI2XL U1720 ( .A(n1604), .B(n3599), .S0(n331), .Y(n2844) );
  MXI2XL U1721 ( .A(n1605), .B(n3598), .S0(n332), .Y(n2845) );
  MXI2XL U1722 ( .A(n1606), .B(n3597), .S0(n335), .Y(n2846) );
  MXI2XL U1723 ( .A(n1607), .B(n3596), .S0(n339), .Y(n2847) );
  MXI2XL U1724 ( .A(n1608), .B(n3595), .S0(n336), .Y(n2848) );
  MXI2XL U1725 ( .A(n1609), .B(n3594), .S0(n334), .Y(n2849) );
  MXI2XL U1726 ( .A(n1610), .B(n3593), .S0(n338), .Y(n2850) );
  MXI2XL U1727 ( .A(n1611), .B(n3592), .S0(n331), .Y(n2851) );
  MXI2XL U1728 ( .A(n1612), .B(n3591), .S0(n332), .Y(n2852) );
  MXI2XL U1729 ( .A(n1613), .B(n3590), .S0(n335), .Y(n2853) );
  MXI2XL U1730 ( .A(n1614), .B(n3589), .S0(n339), .Y(n2854) );
  MXI2XL U1731 ( .A(n1615), .B(n3588), .S0(n339), .Y(n2855) );
  MXI2XL U1732 ( .A(n1616), .B(n3587), .S0(n339), .Y(n2856) );
  MXI2XL U1733 ( .A(n1617), .B(n3586), .S0(n339), .Y(n2857) );
  MXI2XL U1734 ( .A(n1618), .B(n3585), .S0(n339), .Y(n2858) );
  MXI2XL U1735 ( .A(n1619), .B(n3584), .S0(n339), .Y(n2859) );
  MXI2XL U1736 ( .A(n1620), .B(n3583), .S0(n339), .Y(n2860) );
  MXI2XL U1737 ( .A(n1621), .B(n3582), .S0(n339), .Y(n2861) );
  MXI2XL U1738 ( .A(n1622), .B(n3581), .S0(n339), .Y(n2862) );
  MXI2XL U1739 ( .A(n1623), .B(n3580), .S0(n339), .Y(n2863) );
  MXI2XL U1740 ( .A(n1754), .B(n3604), .S0(n326), .Y(n2994) );
  MXI2XL U1741 ( .A(n1755), .B(n3603), .S0(n330), .Y(n2995) );
  MXI2XL U1742 ( .A(n1756), .B(n3602), .S0(n327), .Y(n2996) );
  MXI2XL U1743 ( .A(n1757), .B(n3601), .S0(n325), .Y(n2997) );
  MXI2XL U1744 ( .A(n1758), .B(n3600), .S0(n329), .Y(n2998) );
  MXI2XL U1745 ( .A(n1759), .B(n3599), .S0(n322), .Y(n2999) );
  MXI2XL U1746 ( .A(n1760), .B(n3598), .S0(n323), .Y(n3000) );
  MXI2XL U1747 ( .A(n1761), .B(n3597), .S0(n326), .Y(n3001) );
  MXI2XL U1748 ( .A(n1762), .B(n3596), .S0(n330), .Y(n3002) );
  MXI2XL U1749 ( .A(n1763), .B(n3595), .S0(n327), .Y(n3003) );
  MXI2XL U1750 ( .A(n1764), .B(n3594), .S0(n325), .Y(n3004) );
  MXI2XL U1751 ( .A(n1765), .B(n3593), .S0(n329), .Y(n3005) );
  MXI2XL U1752 ( .A(n1766), .B(n3592), .S0(n322), .Y(n3006) );
  MXI2XL U1753 ( .A(n1767), .B(n3591), .S0(n323), .Y(n3007) );
  MXI2XL U1754 ( .A(n1768), .B(n3590), .S0(n326), .Y(n3008) );
  MXI2XL U1755 ( .A(n1769), .B(n3589), .S0(n330), .Y(n3009) );
  MXI2XL U1756 ( .A(n1770), .B(n3588), .S0(n330), .Y(n3010) );
  MXI2XL U1757 ( .A(n1771), .B(n3587), .S0(n330), .Y(n3011) );
  MXI2XL U1758 ( .A(n1772), .B(n3586), .S0(n330), .Y(n3012) );
  MXI2XL U1759 ( .A(n1773), .B(n3585), .S0(n330), .Y(n3013) );
  MXI2XL U1760 ( .A(n1774), .B(n3584), .S0(n330), .Y(n3014) );
  MXI2XL U1761 ( .A(n1775), .B(n3583), .S0(n330), .Y(n3015) );
  MXI2XL U1762 ( .A(n1776), .B(n3582), .S0(n330), .Y(n3016) );
  MXI2XL U1763 ( .A(n1777), .B(n3581), .S0(n330), .Y(n3017) );
  MXI2XL U1764 ( .A(n1778), .B(n3580), .S0(n330), .Y(n3018) );
  XOR2XL U1765 ( .A(proc_addr[7]), .B(N57), .Y(n3800) );
  XOR2XL U1766 ( .A(proc_addr[6]), .B(N58), .Y(n3798) );
  MXI2XL U1767 ( .A(n695), .B(n3577), .S0(n393), .Y(n1935) );
  MXI2XL U1768 ( .A(n850), .B(n3577), .S0(n384), .Y(n2090) );
  MXI2XL U1769 ( .A(n1005), .B(n3577), .S0(n375), .Y(n2245) );
  MXI2XL U1770 ( .A(n1160), .B(n3577), .S0(n366), .Y(n2400) );
  MXI2XL U1771 ( .A(n1315), .B(n3577), .S0(n357), .Y(n2555) );
  MXI2XL U1772 ( .A(n1470), .B(n3577), .S0(n348), .Y(n2710) );
  MXI2XL U1773 ( .A(n1625), .B(n3577), .S0(n339), .Y(n2865) );
  MXI2XL U1774 ( .A(n1780), .B(n3577), .S0(n330), .Y(n3021) );
  MXI2XL U1775 ( .A(n694), .B(n3579), .S0(n393), .Y(n1934) );
  MXI2XL U1776 ( .A(n849), .B(n3579), .S0(n384), .Y(n2089) );
  MXI2XL U1777 ( .A(n1004), .B(n3579), .S0(n375), .Y(n2244) );
  MXI2XL U1778 ( .A(n1159), .B(n3579), .S0(n366), .Y(n2399) );
  MXI2XL U1779 ( .A(n1314), .B(n3579), .S0(n357), .Y(n2554) );
  MXI2XL U1780 ( .A(n1469), .B(n3579), .S0(n348), .Y(n2709) );
  MXI2XL U1781 ( .A(n1624), .B(n3579), .S0(n339), .Y(n2864) );
  MXI2XL U1782 ( .A(n1779), .B(n3579), .S0(n330), .Y(n3019) );
  XNOR2XL U1783 ( .A(N35), .B(proc_addr[29]), .Y(n3782) );
  XNOR2XL U1784 ( .A(N37), .B(proc_addr[27]), .Y(n3780) );
  XNOR2XL U1785 ( .A(N36), .B(proc_addr[28]), .Y(n3781) );
  XNOR2XL U1786 ( .A(N43), .B(proc_addr[21]), .Y(n3789) );
  XNOR2XL U1787 ( .A(N44), .B(proc_addr[20]), .Y(n3788) );
  XNOR2XL U1788 ( .A(N42), .B(proc_addr[22]), .Y(n3787) );
  XNOR2XL U1789 ( .A(N49), .B(proc_addr[15]), .Y(n3796) );
  XNOR2XL U1790 ( .A(N50), .B(proc_addr[14]), .Y(n3795) );
  XNOR2XL U1791 ( .A(N48), .B(proc_addr[16]), .Y(n3794) );
  CLKINVX1 U1792 ( .A(N32), .Y(n475) );
  CLKINVX1 U1793 ( .A(N30), .Y(n439) );
  CLKINVX1 U1794 ( .A(N31), .Y(n463) );
  CLKBUFX3 U1795 ( .A(n393), .Y(n385) );
  CLKBUFX3 U1796 ( .A(n393), .Y(n386) );
  CLKBUFX3 U1797 ( .A(n393), .Y(n387) );
  CLKBUFX3 U1798 ( .A(n390), .Y(n388) );
  CLKBUFX3 U1799 ( .A(n393), .Y(n389) );
  CLKBUFX3 U1800 ( .A(n3739), .Y(n390) );
  CLKBUFX3 U1801 ( .A(n390), .Y(n391) );
  CLKBUFX3 U1802 ( .A(n390), .Y(n392) );
  CLKBUFX3 U1803 ( .A(n384), .Y(n376) );
  CLKBUFX3 U1804 ( .A(n384), .Y(n377) );
  CLKBUFX3 U1805 ( .A(n384), .Y(n378) );
  CLKBUFX3 U1806 ( .A(n381), .Y(n379) );
  CLKBUFX3 U1807 ( .A(n384), .Y(n380) );
  CLKBUFX3 U1808 ( .A(n3738), .Y(n381) );
  CLKBUFX3 U1809 ( .A(n381), .Y(n382) );
  CLKBUFX3 U1810 ( .A(n381), .Y(n383) );
  CLKBUFX3 U1811 ( .A(n375), .Y(n367) );
  CLKBUFX3 U1812 ( .A(n375), .Y(n368) );
  CLKBUFX3 U1813 ( .A(n375), .Y(n369) );
  CLKBUFX3 U1814 ( .A(n372), .Y(n370) );
  CLKBUFX3 U1815 ( .A(n375), .Y(n371) );
  CLKBUFX3 U1816 ( .A(n3737), .Y(n372) );
  CLKBUFX3 U1817 ( .A(n372), .Y(n373) );
  CLKBUFX3 U1818 ( .A(n372), .Y(n374) );
  CLKBUFX3 U1819 ( .A(n366), .Y(n358) );
  CLKBUFX3 U1820 ( .A(n366), .Y(n359) );
  CLKBUFX3 U1821 ( .A(n366), .Y(n360) );
  CLKBUFX3 U1822 ( .A(n363), .Y(n361) );
  CLKBUFX3 U1823 ( .A(n366), .Y(n362) );
  CLKBUFX3 U1824 ( .A(n3736), .Y(n363) );
  CLKBUFX3 U1825 ( .A(n363), .Y(n364) );
  CLKBUFX3 U1826 ( .A(n363), .Y(n365) );
  CLKBUFX3 U1827 ( .A(n3739), .Y(n393) );
  CLKBUFX3 U1828 ( .A(n3738), .Y(n384) );
  CLKBUFX3 U1829 ( .A(n3737), .Y(n375) );
  CLKBUFX3 U1830 ( .A(n3736), .Y(n366) );
  CLKBUFX3 U1831 ( .A(n357), .Y(n349) );
  CLKBUFX3 U1832 ( .A(n357), .Y(n350) );
  CLKBUFX3 U1833 ( .A(n357), .Y(n351) );
  CLKBUFX3 U1834 ( .A(n354), .Y(n352) );
  CLKBUFX3 U1835 ( .A(n357), .Y(n353) );
  CLKBUFX3 U1836 ( .A(n3735), .Y(n354) );
  CLKBUFX3 U1837 ( .A(n354), .Y(n355) );
  CLKBUFX3 U1838 ( .A(n354), .Y(n356) );
  CLKBUFX3 U1839 ( .A(n348), .Y(n340) );
  CLKBUFX3 U1840 ( .A(n348), .Y(n341) );
  CLKBUFX3 U1841 ( .A(n348), .Y(n342) );
  CLKBUFX3 U1842 ( .A(n345), .Y(n343) );
  CLKBUFX3 U1843 ( .A(n348), .Y(n344) );
  CLKBUFX3 U1844 ( .A(n3734), .Y(n345) );
  CLKBUFX3 U1845 ( .A(n345), .Y(n346) );
  CLKBUFX3 U1846 ( .A(n345), .Y(n347) );
  CLKBUFX3 U1847 ( .A(n339), .Y(n331) );
  CLKBUFX3 U1848 ( .A(n339), .Y(n332) );
  CLKBUFX3 U1849 ( .A(n339), .Y(n333) );
  CLKBUFX3 U1850 ( .A(n336), .Y(n334) );
  CLKBUFX3 U1851 ( .A(n339), .Y(n335) );
  CLKBUFX3 U1852 ( .A(n3733), .Y(n336) );
  CLKBUFX3 U1853 ( .A(n336), .Y(n337) );
  CLKBUFX3 U1854 ( .A(n336), .Y(n338) );
  CLKBUFX3 U1855 ( .A(n330), .Y(n322) );
  CLKBUFX3 U1856 ( .A(n330), .Y(n323) );
  CLKBUFX3 U1857 ( .A(n330), .Y(n324) );
  CLKBUFX3 U1858 ( .A(n327), .Y(n325) );
  CLKBUFX3 U1859 ( .A(n330), .Y(n326) );
  CLKBUFX3 U1860 ( .A(n3578), .Y(n327) );
  CLKBUFX3 U1861 ( .A(n327), .Y(n328) );
  CLKBUFX3 U1862 ( .A(n327), .Y(n329) );
  CLKBUFX3 U1863 ( .A(n3735), .Y(n357) );
  CLKBUFX3 U1864 ( .A(n3734), .Y(n348) );
  CLKBUFX3 U1865 ( .A(n3733), .Y(n339) );
  CLKBUFX3 U1866 ( .A(n3578), .Y(n330) );
  CLKBUFX3 U1867 ( .A(n3065), .Y(n3039) );
  CLKBUFX3 U1868 ( .A(n3068), .Y(n3025) );
  CLKBUFX3 U1869 ( .A(n3070), .Y(n537) );
  CLKBUFX3 U1870 ( .A(n3072), .Y(n529) );
  CLKBUFX3 U1871 ( .A(n3074), .Y(n521) );
  CLKBUFX3 U1872 ( .A(n3076), .Y(n513) );
  CLKBUFX3 U1873 ( .A(n3060), .Y(n3058) );
  CLKBUFX3 U1874 ( .A(n3078), .Y(n505) );
  CLKBUFX3 U1875 ( .A(n3080), .Y(n497) );
  CLKBUFX3 U1876 ( .A(n3082), .Y(n489) );
  CLKBUFX3 U1877 ( .A(n3067), .Y(n3031) );
  CLKBUFX3 U1878 ( .A(n3067), .Y(n3028) );
  CLKBUFX3 U1879 ( .A(n3065), .Y(n3038) );
  CLKBUFX3 U1880 ( .A(n3069), .Y(n3023) );
  CLKBUFX3 U1881 ( .A(n3069), .Y(n540) );
  CLKBUFX3 U1882 ( .A(n3071), .Y(n535) );
  CLKBUFX3 U1883 ( .A(n3071), .Y(n532) );
  CLKBUFX3 U1884 ( .A(n3073), .Y(n527) );
  CLKBUFX3 U1885 ( .A(n3073), .Y(n524) );
  CLKBUFX3 U1886 ( .A(n3075), .Y(n519) );
  CLKBUFX3 U1887 ( .A(n3075), .Y(n516) );
  CLKBUFX3 U1888 ( .A(n3077), .Y(n511) );
  CLKBUFX3 U1889 ( .A(n3065), .Y(n3037) );
  CLKBUFX3 U1890 ( .A(n3077), .Y(n508) );
  CLKBUFX3 U1891 ( .A(n3079), .Y(n503) );
  CLKBUFX3 U1892 ( .A(n3079), .Y(n500) );
  CLKBUFX3 U1893 ( .A(n3081), .Y(n495) );
  CLKBUFX3 U1894 ( .A(n3081), .Y(n492) );
  CLKBUFX3 U1895 ( .A(n3083), .Y(n487) );
  CLKBUFX3 U1896 ( .A(n3083), .Y(n484) );
  CLKBUFX3 U1897 ( .A(n3067), .Y(n3029) );
  CLKBUFX3 U1898 ( .A(n3068), .Y(n3026) );
  CLKBUFX3 U1899 ( .A(n3065), .Y(n3036) );
  CLKBUFX3 U1900 ( .A(n3069), .Y(n3020) );
  CLKBUFX3 U1901 ( .A(n3070), .Y(n538) );
  CLKBUFX3 U1902 ( .A(n3071), .Y(n533) );
  CLKBUFX3 U1903 ( .A(n3072), .Y(n530) );
  CLKBUFX3 U1904 ( .A(n3073), .Y(n525) );
  CLKBUFX3 U1905 ( .A(n3074), .Y(n522) );
  CLKBUFX3 U1906 ( .A(n3075), .Y(n517) );
  CLKBUFX3 U1907 ( .A(n3076), .Y(n514) );
  CLKBUFX3 U1908 ( .A(n3066), .Y(n3035) );
  CLKBUFX3 U1909 ( .A(n3077), .Y(n509) );
  CLKBUFX3 U1910 ( .A(n3078), .Y(n506) );
  CLKBUFX3 U1911 ( .A(n3079), .Y(n501) );
  CLKBUFX3 U1912 ( .A(n3080), .Y(n498) );
  CLKBUFX3 U1913 ( .A(n3081), .Y(n493) );
  CLKBUFX3 U1914 ( .A(n3082), .Y(n490) );
  CLKBUFX3 U1915 ( .A(n3083), .Y(n485) );
  CLKBUFX3 U1916 ( .A(n3066), .Y(n3032) );
  CLKBUFX3 U1917 ( .A(n3067), .Y(n3030) );
  CLKBUFX3 U1918 ( .A(n3068), .Y(n3027) );
  CLKBUFX3 U1919 ( .A(n3066), .Y(n3034) );
  CLKBUFX3 U1920 ( .A(n3068), .Y(n3024) );
  CLKBUFX3 U1921 ( .A(n3069), .Y(n3022) );
  CLKBUFX3 U1922 ( .A(n3070), .Y(n539) );
  CLKBUFX3 U1923 ( .A(n3070), .Y(n536) );
  CLKBUFX3 U1924 ( .A(n3071), .Y(n534) );
  CLKBUFX3 U1925 ( .A(n3072), .Y(n531) );
  CLKBUFX3 U1926 ( .A(n3072), .Y(n528) );
  CLKBUFX3 U1927 ( .A(n3073), .Y(n526) );
  CLKBUFX3 U1928 ( .A(n3074), .Y(n523) );
  CLKBUFX3 U1929 ( .A(n3074), .Y(n520) );
  CLKBUFX3 U1930 ( .A(n3075), .Y(n518) );
  CLKBUFX3 U1931 ( .A(n3076), .Y(n515) );
  CLKBUFX3 U1932 ( .A(n3076), .Y(n512) );
  CLKBUFX3 U1933 ( .A(n3066), .Y(n3033) );
  CLKBUFX3 U1934 ( .A(n3077), .Y(n510) );
  CLKBUFX3 U1935 ( .A(n3078), .Y(n507) );
  CLKBUFX3 U1936 ( .A(n3078), .Y(n504) );
  CLKBUFX3 U1937 ( .A(n3079), .Y(n502) );
  CLKBUFX3 U1938 ( .A(n3080), .Y(n499) );
  CLKBUFX3 U1939 ( .A(n3080), .Y(n496) );
  CLKBUFX3 U1940 ( .A(n3081), .Y(n494) );
  CLKBUFX3 U1941 ( .A(n3082), .Y(n491) );
  CLKBUFX3 U1942 ( .A(n3082), .Y(n488) );
  CLKBUFX3 U1943 ( .A(n3083), .Y(n486) );
  CLKBUFX3 U1944 ( .A(n3061), .Y(n3055) );
  CLKBUFX3 U1945 ( .A(n3061), .Y(n3054) );
  CLKBUFX3 U1946 ( .A(n3061), .Y(n3053) );
  CLKBUFX3 U1947 ( .A(n3061), .Y(n3052) );
  CLKBUFX3 U1948 ( .A(n3062), .Y(n3051) );
  CLKBUFX3 U1949 ( .A(n3062), .Y(n3050) );
  CLKBUFX3 U1950 ( .A(n3062), .Y(n3049) );
  CLKBUFX3 U1951 ( .A(n3062), .Y(n3048) );
  CLKBUFX3 U1952 ( .A(n3063), .Y(n3047) );
  CLKBUFX3 U1953 ( .A(n3063), .Y(n3046) );
  CLKBUFX3 U1954 ( .A(n3063), .Y(n3045) );
  CLKBUFX3 U1955 ( .A(n3063), .Y(n3044) );
  CLKBUFX3 U1956 ( .A(n3064), .Y(n3043) );
  CLKBUFX3 U1957 ( .A(n3064), .Y(n3042) );
  CLKBUFX3 U1958 ( .A(n3064), .Y(n3041) );
  CLKBUFX3 U1959 ( .A(n3064), .Y(n3040) );
  CLKBUFX3 U1960 ( .A(n3060), .Y(n3056) );
  CLKBUFX3 U1961 ( .A(n3060), .Y(n3057) );
  INVX3 U1962 ( .A(n413), .Y(n405) );
  INVX3 U1963 ( .A(n417), .Y(n406) );
  INVX3 U1964 ( .A(n417), .Y(n407) );
  INVX3 U1965 ( .A(n417), .Y(n408) );
  INVX3 U1966 ( .A(n319), .Y(n409) );
  INVX3 U1967 ( .A(n416), .Y(n410) );
  INVX3 U1968 ( .A(n413), .Y(n402) );
  INVX3 U1969 ( .A(n416), .Y(n403) );
  INVX3 U1970 ( .A(n416), .Y(n404) );
  INVX3 U1971 ( .A(n319), .Y(n411) );
  CLKBUFX3 U1972 ( .A(n3060), .Y(n3059) );
  INVX3 U1973 ( .A(n417), .Y(n412) );
  INVX3 U1974 ( .A(n438), .Y(n426) );
  INVX3 U1975 ( .A(n437), .Y(n427) );
  INVX3 U1976 ( .A(n437), .Y(n428) );
  INVX3 U1977 ( .A(n438), .Y(n429) );
  INVX3 U1978 ( .A(n437), .Y(n430) );
  INVX3 U1979 ( .A(n437), .Y(n431) );
  INVX3 U1980 ( .A(n439), .Y(n432) );
  INVX3 U1981 ( .A(n439), .Y(n433) );
  INVX3 U1982 ( .A(n437), .Y(n434) );
  INVX3 U1983 ( .A(n437), .Y(n435) );
  INVX3 U1984 ( .A(n437), .Y(n418) );
  INVX3 U1985 ( .A(n437), .Y(n419) );
  INVX3 U1986 ( .A(n437), .Y(n420) );
  INVX3 U1987 ( .A(n438), .Y(n421) );
  INVX3 U1988 ( .A(n437), .Y(n422) );
  INVX3 U1989 ( .A(n438), .Y(n423) );
  INVX3 U1990 ( .A(n438), .Y(n424) );
  INVX3 U1991 ( .A(n438), .Y(n425) );
  CLKBUFX3 U1992 ( .A(n3084), .Y(n481) );
  CLKBUFX3 U1993 ( .A(n3085), .Y(n479) );
  CLKBUFX3 U1994 ( .A(n3085), .Y(n476) );
  CLKBUFX3 U1995 ( .A(n3084), .Y(n482) );
  CLKBUFX3 U1996 ( .A(n3085), .Y(n477) );
  CLKBUFX3 U1997 ( .A(n3084), .Y(n483) );
  CLKBUFX3 U1998 ( .A(n3084), .Y(n480) );
  CLKBUFX3 U1999 ( .A(n3085), .Y(n478) );
  INVX3 U2000 ( .A(n461), .Y(n460) );
  CLKBUFX3 U2001 ( .A(n413), .Y(n415) );
  INVX3 U2002 ( .A(n462), .Y(n440) );
  INVX3 U2003 ( .A(n461), .Y(n441) );
  INVX3 U2004 ( .A(n462), .Y(n442) );
  INVX3 U2005 ( .A(n461), .Y(n443) );
  INVX3 U2006 ( .A(n461), .Y(n444) );
  INVX3 U2007 ( .A(n462), .Y(n445) );
  INVX3 U2008 ( .A(n461), .Y(n446) );
  INVX3 U2009 ( .A(n462), .Y(n447) );
  INVX3 U2010 ( .A(n462), .Y(n448) );
  INVX3 U2011 ( .A(n462), .Y(n449) );
  INVX3 U2012 ( .A(n462), .Y(n450) );
  CLKBUFX3 U2013 ( .A(n416), .Y(n413) );
  INVX3 U2014 ( .A(n462), .Y(n451) );
  INVX3 U2015 ( .A(n462), .Y(n452) );
  INVX3 U2016 ( .A(n463), .Y(n453) );
  INVX3 U2017 ( .A(n463), .Y(n454) );
  INVX3 U2018 ( .A(n461), .Y(n455) );
  INVX3 U2019 ( .A(n462), .Y(n456) );
  INVX3 U2020 ( .A(n461), .Y(n457) );
  INVX3 U2021 ( .A(n461), .Y(n458) );
  INVX3 U2022 ( .A(n461), .Y(n459) );
  CLKBUFX3 U2023 ( .A(n319), .Y(mem_write) );
  CLKBUFX3 U2024 ( .A(n3093), .Y(n3065) );
  CLKBUFX3 U2025 ( .A(n3090), .Y(n3067) );
  CLKBUFX3 U2026 ( .A(n3089), .Y(n3068) );
  CLKBUFX3 U2027 ( .A(n3089), .Y(n3069) );
  CLKBUFX3 U2028 ( .A(n3094), .Y(n3070) );
  CLKBUFX3 U2029 ( .A(n3094), .Y(n3071) );
  CLKBUFX3 U2030 ( .A(n3088), .Y(n3072) );
  CLKBUFX3 U2031 ( .A(n3088), .Y(n3073) );
  CLKBUFX3 U2032 ( .A(n3095), .Y(n3074) );
  CLKBUFX3 U2033 ( .A(n3095), .Y(n3075) );
  CLKBUFX3 U2034 ( .A(n3087), .Y(n3076) );
  CLKBUFX3 U2035 ( .A(n3090), .Y(n3066) );
  CLKBUFX3 U2036 ( .A(n3087), .Y(n3077) );
  CLKBUFX3 U2037 ( .A(n3096), .Y(n3078) );
  CLKBUFX3 U2038 ( .A(n3096), .Y(n3079) );
  CLKBUFX3 U2039 ( .A(n3086), .Y(n3080) );
  CLKBUFX3 U2040 ( .A(n3086), .Y(n3081) );
  CLKBUFX3 U2041 ( .A(n3097), .Y(n3082) );
  CLKBUFX3 U2042 ( .A(n3097), .Y(n3083) );
  CLKBUFX3 U2043 ( .A(n3092), .Y(n3061) );
  CLKBUFX3 U2044 ( .A(n3091), .Y(n3062) );
  CLKBUFX3 U2045 ( .A(n3091), .Y(n3063) );
  CLKBUFX3 U2046 ( .A(n3089), .Y(n3064) );
  CLKBUFX3 U2047 ( .A(n3092), .Y(n3060) );
  INVX3 U2048 ( .A(n438), .Y(n436) );
  INVX3 U2049 ( .A(n475), .Y(n472) );
  INVX3 U2050 ( .A(n474), .Y(n464) );
  INVX3 U2051 ( .A(n474), .Y(n465) );
  INVX3 U2052 ( .A(n474), .Y(n466) );
  INVX3 U2053 ( .A(n474), .Y(n467) );
  INVX3 U2054 ( .A(n474), .Y(n468) );
  INVX3 U2055 ( .A(n474), .Y(n469) );
  INVX3 U2056 ( .A(n474), .Y(n470) );
  INVX3 U2057 ( .A(n475), .Y(n471) );
  CLKBUFX3 U2058 ( .A(n439), .Y(n437) );
  CLKBUFX3 U2059 ( .A(n462), .Y(n461) );
  CLKBUFX3 U2060 ( .A(n439), .Y(n438) );
  CLKBUFX3 U2061 ( .A(n463), .Y(n462) );
  CLKBUFX3 U2062 ( .A(n401), .Y(n400) );
  CLKBUFX3 U2063 ( .A(n3744), .Y(n399) );
  CLKBUFX3 U2064 ( .A(n399), .Y(n398) );
  CLKBUFX3 U2065 ( .A(n396), .Y(n397) );
  CLKBUFX3 U2066 ( .A(n3744), .Y(n396) );
  CLKBUFX3 U2067 ( .A(n396), .Y(n395) );
  CLKBUFX3 U2068 ( .A(n3744), .Y(n401) );
  CLKBUFX3 U2069 ( .A(n3744), .Y(n394) );
  CLKBUFX3 U2070 ( .A(n319), .Y(n416) );
  CLKBUFX3 U2071 ( .A(n3094), .Y(n3089) );
  CLKBUFX3 U2072 ( .A(n3095), .Y(n3088) );
  CLKBUFX3 U2073 ( .A(n3096), .Y(n3087) );
  CLKBUFX3 U2074 ( .A(n3097), .Y(n3086) );
  CLKBUFX3 U2075 ( .A(n3093), .Y(n3090) );
  CLKBUFX3 U2076 ( .A(n3092), .Y(n3091) );
  CLKBUFX3 U2077 ( .A(n3099), .Y(n3084) );
  CLKBUFX3 U2078 ( .A(n3093), .Y(n3085) );
  CLKINVX1 U2079 ( .A(n474), .Y(n473) );
  CLKBUFX3 U2080 ( .A(n475), .Y(n474) );
  CLKBUFX3 U2081 ( .A(n3098), .Y(n3094) );
  CLKBUFX3 U2082 ( .A(n3098), .Y(n3095) );
  CLKBUFX3 U2083 ( .A(n3098), .Y(n3096) );
  CLKBUFX2 U2084 ( .A(n3098), .Y(n3097) );
  CLKBUFX3 U2085 ( .A(n3099), .Y(n3093) );
  CLKBUFX3 U2086 ( .A(n3099), .Y(n3092) );
  CLKBUFX3 U2087 ( .A(n319), .Y(n417) );
  CLKINVX1 U2088 ( .A(proc_reset), .Y(n3098) );
  INVXL U2089 ( .A(proc_reset), .Y(n3099) );
  AND4X1 U2090 ( .A(N34), .B(n3770), .C(n3763), .D(n3743), .Y(n319) );
  CLKMX2X2 U2091 ( .A(n320), .B(n321), .S0(n472), .Y(N34) );
  MX4X1 U2092 ( .A(\CACHE[0][153] ), .B(\CACHE[1][153] ), .C(\CACHE[2][153] ), 
        .D(\CACHE[3][153] ), .S0(n421), .S1(n460), .Y(n320) );
  MX4X1 U2093 ( .A(\CACHE[4][153] ), .B(\CACHE[5][153] ), .C(\CACHE[6][153] ), 
        .D(\CACHE[7][153] ), .S0(n436), .S1(n460), .Y(n321) );
  MXI2X1 U2094 ( .A(n3362), .B(n3363), .S0(n466), .Y(N56) );
  MXI4X1 U2095 ( .A(\CACHE[4][131] ), .B(\CACHE[5][131] ), .C(\CACHE[6][131] ), 
        .D(\CACHE[7][131] ), .S0(n423), .S1(n457), .Y(n3363) );
  MXI4X1 U2096 ( .A(\CACHE[0][131] ), .B(\CACHE[1][131] ), .C(\CACHE[2][131] ), 
        .D(\CACHE[3][131] ), .S0(n423), .S1(n457), .Y(n3362) );
  MXI2X1 U2097 ( .A(n3364), .B(n3365), .S0(n471), .Y(N55) );
  MXI4X1 U2098 ( .A(\CACHE[4][132] ), .B(\CACHE[5][132] ), .C(\CACHE[6][132] ), 
        .D(\CACHE[7][132] ), .S0(n423), .S1(n442), .Y(n3365) );
  MXI4X1 U2099 ( .A(\CACHE[0][132] ), .B(\CACHE[1][132] ), .C(\CACHE[2][132] ), 
        .D(\CACHE[3][132] ), .S0(n423), .S1(n440), .Y(n3364) );
  MXI2X1 U2100 ( .A(n3366), .B(n3367), .S0(n471), .Y(N54) );
  MXI4X1 U2101 ( .A(\CACHE[4][133] ), .B(\CACHE[5][133] ), .C(\CACHE[6][133] ), 
        .D(\CACHE[7][133] ), .S0(n423), .S1(n451), .Y(n3367) );
  MXI4X1 U2102 ( .A(\CACHE[0][133] ), .B(\CACHE[1][133] ), .C(\CACHE[2][133] ), 
        .D(\CACHE[3][133] ), .S0(n423), .S1(n450), .Y(n3366) );
  MXI2X1 U2103 ( .A(n3374), .B(n3375), .S0(n471), .Y(N50) );
  MXI4X1 U2104 ( .A(\CACHE[4][137] ), .B(\CACHE[5][137] ), .C(\CACHE[6][137] ), 
        .D(\CACHE[7][137] ), .S0(n424), .S1(n441), .Y(n3375) );
  MXI4X1 U2105 ( .A(\CACHE[0][137] ), .B(\CACHE[1][137] ), .C(\CACHE[2][137] ), 
        .D(\CACHE[3][137] ), .S0(n424), .S1(n458), .Y(n3374) );
  MXI2X1 U2106 ( .A(n3376), .B(n3377), .S0(n471), .Y(N49) );
  MXI4X1 U2107 ( .A(\CACHE[4][138] ), .B(\CACHE[5][138] ), .C(\CACHE[6][138] ), 
        .D(\CACHE[7][138] ), .S0(n424), .S1(n458), .Y(n3377) );
  MXI4X1 U2108 ( .A(\CACHE[0][138] ), .B(\CACHE[1][138] ), .C(\CACHE[2][138] ), 
        .D(\CACHE[3][138] ), .S0(n424), .S1(n458), .Y(n3376) );
  MXI2X1 U2109 ( .A(n3378), .B(n3379), .S0(n471), .Y(N48) );
  MXI4X1 U2110 ( .A(\CACHE[4][139] ), .B(\CACHE[5][139] ), .C(\CACHE[6][139] ), 
        .D(\CACHE[7][139] ), .S0(n424), .S1(n458), .Y(n3379) );
  MXI4X1 U2111 ( .A(\CACHE[0][139] ), .B(\CACHE[1][139] ), .C(\CACHE[2][139] ), 
        .D(\CACHE[3][139] ), .S0(n424), .S1(n458), .Y(n3378) );
  MXI2X1 U2112 ( .A(n3386), .B(n3387), .S0(n471), .Y(N44) );
  MXI4X1 U2113 ( .A(\CACHE[4][143] ), .B(\CACHE[5][143] ), .C(\CACHE[6][143] ), 
        .D(\CACHE[7][143] ), .S0(n425), .S1(n458), .Y(n3387) );
  MXI4X1 U2114 ( .A(\CACHE[0][143] ), .B(\CACHE[1][143] ), .C(\CACHE[2][143] ), 
        .D(\CACHE[3][143] ), .S0(n425), .S1(n458), .Y(n3386) );
  MXI2X1 U2115 ( .A(n3388), .B(n3389), .S0(n472), .Y(N43) );
  MXI4X1 U2116 ( .A(\CACHE[4][144] ), .B(\CACHE[5][144] ), .C(\CACHE[6][144] ), 
        .D(\CACHE[7][144] ), .S0(n425), .S1(n459), .Y(n3389) );
  MXI4X1 U2117 ( .A(\CACHE[0][144] ), .B(\CACHE[1][144] ), .C(\CACHE[2][144] ), 
        .D(\CACHE[3][144] ), .S0(n425), .S1(n459), .Y(n3388) );
  MXI2X1 U2118 ( .A(n3390), .B(n3391), .S0(n472), .Y(N42) );
  MXI4X1 U2119 ( .A(\CACHE[4][145] ), .B(\CACHE[5][145] ), .C(\CACHE[6][145] ), 
        .D(\CACHE[7][145] ), .S0(n425), .S1(n459), .Y(n3391) );
  MXI4X1 U2120 ( .A(\CACHE[0][145] ), .B(\CACHE[1][145] ), .C(\CACHE[2][145] ), 
        .D(\CACHE[3][145] ), .S0(n425), .S1(n459), .Y(n3390) );
  MXI2X1 U2121 ( .A(n3398), .B(n3399), .S0(n472), .Y(N38) );
  MXI4X1 U2122 ( .A(\CACHE[4][149] ), .B(\CACHE[5][149] ), .C(\CACHE[6][149] ), 
        .D(\CACHE[7][149] ), .S0(n433), .S1(n459), .Y(n3399) );
  MXI4X1 U2123 ( .A(\CACHE[0][149] ), .B(\CACHE[1][149] ), .C(\CACHE[2][149] ), 
        .D(\CACHE[3][149] ), .S0(n432), .S1(n459), .Y(n3398) );
  MXI2X1 U2124 ( .A(n3400), .B(n3401), .S0(n472), .Y(N37) );
  MXI4X1 U2125 ( .A(\CACHE[4][150] ), .B(\CACHE[5][150] ), .C(\CACHE[6][150] ), 
        .D(\CACHE[7][150] ), .S0(n430), .S1(n460), .Y(n3401) );
  MXI4X1 U2126 ( .A(\CACHE[0][150] ), .B(\CACHE[1][150] ), .C(\CACHE[2][150] ), 
        .D(\CACHE[3][150] ), .S0(n427), .S1(n460), .Y(n3400) );
  MXI2X1 U2127 ( .A(n3402), .B(n3403), .S0(n472), .Y(N36) );
  MXI4X1 U2128 ( .A(\CACHE[4][151] ), .B(\CACHE[5][151] ), .C(\CACHE[6][151] ), 
        .D(\CACHE[7][151] ), .S0(n435), .S1(n460), .Y(n3403) );
  MXI4X1 U2129 ( .A(\CACHE[0][151] ), .B(\CACHE[1][151] ), .C(\CACHE[2][151] ), 
        .D(\CACHE[3][151] ), .S0(n422), .S1(n460), .Y(n3402) );
  MXI2X1 U2130 ( .A(n3404), .B(n3405), .S0(n472), .Y(N35) );
  MXI4X1 U2131 ( .A(\CACHE[4][152] ), .B(\CACHE[5][152] ), .C(\CACHE[6][152] ), 
        .D(\CACHE[7][152] ), .S0(n420), .S1(n460), .Y(n3405) );
  MXI4X1 U2132 ( .A(\CACHE[0][152] ), .B(\CACHE[1][152] ), .C(\CACHE[2][152] ), 
        .D(\CACHE[3][152] ), .S0(n428), .S1(n460), .Y(n3404) );
  MXI2X1 U2133 ( .A(n3356), .B(n3357), .S0(n469), .Y(N59) );
  MXI4X1 U2134 ( .A(\CACHE[4][128] ), .B(\CACHE[5][128] ), .C(\CACHE[6][128] ), 
        .D(\CACHE[7][128] ), .S0(n422), .S1(n457), .Y(n3357) );
  MXI4X1 U2135 ( .A(\CACHE[0][128] ), .B(\CACHE[1][128] ), .C(\CACHE[2][128] ), 
        .D(\CACHE[3][128] ), .S0(n422), .S1(n457), .Y(n3356) );
  MXI2X1 U2136 ( .A(n3358), .B(n3359), .S0(n470), .Y(N58) );
  MXI4X1 U2137 ( .A(\CACHE[4][129] ), .B(\CACHE[5][129] ), .C(\CACHE[6][129] ), 
        .D(\CACHE[7][129] ), .S0(n422), .S1(n457), .Y(n3359) );
  MXI4X1 U2138 ( .A(\CACHE[0][129] ), .B(\CACHE[1][129] ), .C(\CACHE[2][129] ), 
        .D(\CACHE[3][129] ), .S0(n423), .S1(n457), .Y(n3358) );
  MXI2X1 U2139 ( .A(n3360), .B(n3361), .S0(n472), .Y(N57) );
  MXI4X1 U2140 ( .A(\CACHE[4][130] ), .B(\CACHE[5][130] ), .C(\CACHE[6][130] ), 
        .D(\CACHE[7][130] ), .S0(n423), .S1(n457), .Y(n3361) );
  MXI4X1 U2141 ( .A(\CACHE[0][130] ), .B(\CACHE[1][130] ), .C(\CACHE[2][130] ), 
        .D(\CACHE[3][130] ), .S0(n423), .S1(n457), .Y(n3360) );
  MXI2X1 U2142 ( .A(n3368), .B(n3369), .S0(n471), .Y(N53) );
  MXI4X1 U2143 ( .A(\CACHE[4][134] ), .B(\CACHE[5][134] ), .C(\CACHE[6][134] ), 
        .D(\CACHE[7][134] ), .S0(n423), .S1(n455), .Y(n3369) );
  MXI4X1 U2144 ( .A(\CACHE[0][134] ), .B(\CACHE[1][134] ), .C(\CACHE[2][134] ), 
        .D(\CACHE[3][134] ), .S0(n423), .S1(n446), .Y(n3368) );
  MXI2X1 U2145 ( .A(n3370), .B(n3371), .S0(n471), .Y(N52) );
  MXI4X1 U2146 ( .A(\CACHE[4][135] ), .B(\CACHE[5][135] ), .C(\CACHE[6][135] ), 
        .D(\CACHE[7][135] ), .S0(n423), .S1(n451), .Y(n3371) );
  MXI4X1 U2147 ( .A(\CACHE[0][135] ), .B(\CACHE[1][135] ), .C(\CACHE[2][135] ), 
        .D(\CACHE[3][135] ), .S0(n423), .S1(n457), .Y(n3370) );
  MXI2X1 U2148 ( .A(n3372), .B(n3373), .S0(n471), .Y(N51) );
  MXI4X1 U2149 ( .A(\CACHE[4][136] ), .B(\CACHE[5][136] ), .C(\CACHE[6][136] ), 
        .D(\CACHE[7][136] ), .S0(n424), .S1(n443), .Y(n3373) );
  MXI4X1 U2150 ( .A(\CACHE[0][136] ), .B(\CACHE[1][136] ), .C(\CACHE[2][136] ), 
        .D(\CACHE[3][136] ), .S0(n424), .S1(n459), .Y(n3372) );
  MXI2X1 U2151 ( .A(n3380), .B(n3381), .S0(n471), .Y(N47) );
  MXI4X1 U2152 ( .A(\CACHE[4][140] ), .B(\CACHE[5][140] ), .C(\CACHE[6][140] ), 
        .D(\CACHE[7][140] ), .S0(n424), .S1(n458), .Y(n3381) );
  MXI4X1 U2153 ( .A(\CACHE[0][140] ), .B(\CACHE[1][140] ), .C(\CACHE[2][140] ), 
        .D(\CACHE[3][140] ), .S0(n424), .S1(n458), .Y(n3380) );
  MXI2X1 U2154 ( .A(n3382), .B(n3383), .S0(n471), .Y(N46) );
  MXI4X1 U2155 ( .A(\CACHE[4][141] ), .B(\CACHE[5][141] ), .C(\CACHE[6][141] ), 
        .D(\CACHE[7][141] ), .S0(n424), .S1(n458), .Y(n3383) );
  MXI4X1 U2156 ( .A(\CACHE[0][141] ), .B(\CACHE[1][141] ), .C(\CACHE[2][141] ), 
        .D(\CACHE[3][141] ), .S0(n424), .S1(n458), .Y(n3382) );
  MXI2X1 U2157 ( .A(n3384), .B(n3385), .S0(n471), .Y(N45) );
  MXI4X1 U2158 ( .A(\CACHE[4][142] ), .B(\CACHE[5][142] ), .C(\CACHE[6][142] ), 
        .D(\CACHE[7][142] ), .S0(n424), .S1(n458), .Y(n3385) );
  MXI4X1 U2159 ( .A(\CACHE[0][142] ), .B(\CACHE[1][142] ), .C(\CACHE[2][142] ), 
        .D(\CACHE[3][142] ), .S0(n425), .S1(n458), .Y(n3384) );
  MXI2X1 U2160 ( .A(n3392), .B(n3393), .S0(n472), .Y(N41) );
  MXI4X1 U2161 ( .A(\CACHE[4][146] ), .B(\CACHE[5][146] ), .C(\CACHE[6][146] ), 
        .D(\CACHE[7][146] ), .S0(n425), .S1(n459), .Y(n3393) );
  MXI4X1 U2162 ( .A(\CACHE[0][146] ), .B(\CACHE[1][146] ), .C(\CACHE[2][146] ), 
        .D(\CACHE[3][146] ), .S0(n425), .S1(n459), .Y(n3392) );
  MXI2X1 U2163 ( .A(n3394), .B(n3395), .S0(n472), .Y(N40) );
  MXI4X1 U2164 ( .A(\CACHE[4][147] ), .B(\CACHE[5][147] ), .C(\CACHE[6][147] ), 
        .D(\CACHE[7][147] ), .S0(n425), .S1(n459), .Y(n3395) );
  MXI4X1 U2165 ( .A(\CACHE[0][147] ), .B(\CACHE[1][147] ), .C(\CACHE[2][147] ), 
        .D(\CACHE[3][147] ), .S0(n425), .S1(n459), .Y(n3394) );
  MXI2X1 U2166 ( .A(n3396), .B(n3397), .S0(n472), .Y(N39) );
  MXI4X1 U2167 ( .A(\CACHE[4][148] ), .B(\CACHE[5][148] ), .C(\CACHE[6][148] ), 
        .D(\CACHE[7][148] ), .S0(n425), .S1(n459), .Y(n3397) );
  MXI4X1 U2168 ( .A(\CACHE[0][148] ), .B(\CACHE[1][148] ), .C(\CACHE[2][148] ), 
        .D(\CACHE[3][148] ), .S0(n425), .S1(n459), .Y(n3396) );
  MXI2X1 U2169 ( .A(n3406), .B(n3407), .S0(n472), .Y(N33) );
  MXI4X1 U2170 ( .A(\CACHE[4][154] ), .B(\CACHE[5][154] ), .C(\CACHE[6][154] ), 
        .D(\CACHE[7][154] ), .S0(n431), .S1(n460), .Y(n3407) );
  MXI4X1 U2171 ( .A(\CACHE[0][154] ), .B(\CACHE[1][154] ), .C(\CACHE[2][154] ), 
        .D(\CACHE[3][154] ), .S0(n434), .S1(n460), .Y(n3406) );
  MXI2X1 U2172 ( .A(n3100), .B(n3101), .S0(n464), .Y(N187) );
  MXI4X1 U2173 ( .A(\CACHE[4][0] ), .B(\CACHE[5][0] ), .C(\CACHE[6][0] ), .D(
        \CACHE[7][0] ), .S0(n418), .S1(n440), .Y(n3101) );
  MXI4X1 U2174 ( .A(\CACHE[0][0] ), .B(\CACHE[1][0] ), .C(\CACHE[2][0] ), .D(
        \CACHE[3][0] ), .S0(n430), .S1(n440), .Y(n3100) );
  MXI2X1 U2175 ( .A(n3102), .B(n3103), .S0(n464), .Y(N186) );
  MXI4X1 U2176 ( .A(\CACHE[4][1] ), .B(\CACHE[5][1] ), .C(\CACHE[6][1] ), .D(
        \CACHE[7][1] ), .S0(n426), .S1(n440), .Y(n3103) );
  MXI4X1 U2177 ( .A(\CACHE[0][1] ), .B(\CACHE[1][1] ), .C(\CACHE[2][1] ), .D(
        \CACHE[3][1] ), .S0(n426), .S1(n440), .Y(n3102) );
  MXI2X1 U2178 ( .A(n3104), .B(n3105), .S0(n464), .Y(N185) );
  MXI4X1 U2179 ( .A(\CACHE[4][2] ), .B(\CACHE[5][2] ), .C(\CACHE[6][2] ), .D(
        \CACHE[7][2] ), .S0(n426), .S1(n440), .Y(n3105) );
  MXI4X1 U2180 ( .A(\CACHE[0][2] ), .B(\CACHE[1][2] ), .C(\CACHE[2][2] ), .D(
        \CACHE[3][2] ), .S0(n426), .S1(n440), .Y(n3104) );
  MXI2X1 U2181 ( .A(n3106), .B(n3107), .S0(n464), .Y(N184) );
  MXI4X1 U2182 ( .A(\CACHE[4][3] ), .B(\CACHE[5][3] ), .C(\CACHE[6][3] ), .D(
        \CACHE[7][3] ), .S0(n426), .S1(n440), .Y(n3107) );
  MXI4X1 U2183 ( .A(\CACHE[0][3] ), .B(\CACHE[1][3] ), .C(\CACHE[2][3] ), .D(
        \CACHE[3][3] ), .S0(n426), .S1(n440), .Y(n3106) );
  MXI2X1 U2184 ( .A(n3108), .B(n3109), .S0(n464), .Y(N183) );
  MXI4X1 U2185 ( .A(\CACHE[4][4] ), .B(\CACHE[5][4] ), .C(\CACHE[6][4] ), .D(
        \CACHE[7][4] ), .S0(n426), .S1(n440), .Y(n3109) );
  MXI4X1 U2186 ( .A(\CACHE[0][4] ), .B(\CACHE[1][4] ), .C(\CACHE[2][4] ), .D(
        \CACHE[3][4] ), .S0(n426), .S1(n440), .Y(n3108) );
  MXI2X1 U2187 ( .A(n3110), .B(n3111), .S0(n464), .Y(N182) );
  MXI4X1 U2188 ( .A(\CACHE[4][5] ), .B(\CACHE[5][5] ), .C(\CACHE[6][5] ), .D(
        \CACHE[7][5] ), .S0(n426), .S1(n440), .Y(n3111) );
  MXI4X1 U2189 ( .A(\CACHE[0][5] ), .B(\CACHE[1][5] ), .C(\CACHE[2][5] ), .D(
        \CACHE[3][5] ), .S0(n426), .S1(n440), .Y(n3110) );
  MXI2X1 U2190 ( .A(n3112), .B(n3113), .S0(n464), .Y(N181) );
  MXI4X1 U2191 ( .A(\CACHE[4][6] ), .B(\CACHE[5][6] ), .C(\CACHE[6][6] ), .D(
        \CACHE[7][6] ), .S0(n426), .S1(n441), .Y(n3113) );
  MXI4X1 U2192 ( .A(\CACHE[0][6] ), .B(\CACHE[1][6] ), .C(\CACHE[2][6] ), .D(
        \CACHE[3][6] ), .S0(n426), .S1(n441), .Y(n3112) );
  MXI2X1 U2193 ( .A(n3114), .B(n3115), .S0(n464), .Y(N180) );
  MXI4X1 U2194 ( .A(\CACHE[4][7] ), .B(\CACHE[5][7] ), .C(\CACHE[6][7] ), .D(
        \CACHE[7][7] ), .S0(n426), .S1(n441), .Y(n3115) );
  MXI4X1 U2195 ( .A(\CACHE[0][7] ), .B(\CACHE[1][7] ), .C(\CACHE[2][7] ), .D(
        \CACHE[3][7] ), .S0(n427), .S1(n441), .Y(n3114) );
  MXI2X1 U2196 ( .A(n3116), .B(n3117), .S0(n464), .Y(N179) );
  MXI4X1 U2197 ( .A(\CACHE[4][8] ), .B(\CACHE[5][8] ), .C(\CACHE[6][8] ), .D(
        \CACHE[7][8] ), .S0(n427), .S1(n441), .Y(n3117) );
  MXI4X1 U2198 ( .A(\CACHE[0][8] ), .B(\CACHE[1][8] ), .C(\CACHE[2][8] ), .D(
        \CACHE[3][8] ), .S0(n427), .S1(n441), .Y(n3116) );
  MXI2X1 U2199 ( .A(n3118), .B(n3119), .S0(n464), .Y(N178) );
  MXI4X1 U2200 ( .A(\CACHE[4][9] ), .B(\CACHE[5][9] ), .C(\CACHE[6][9] ), .D(
        \CACHE[7][9] ), .S0(n427), .S1(n441), .Y(n3119) );
  MXI4X1 U2201 ( .A(\CACHE[0][9] ), .B(\CACHE[1][9] ), .C(\CACHE[2][9] ), .D(
        \CACHE[3][9] ), .S0(n427), .S1(n441), .Y(n3118) );
  MXI2X1 U2202 ( .A(n3120), .B(n3121), .S0(n464), .Y(N177) );
  MXI4X1 U2203 ( .A(\CACHE[4][10] ), .B(\CACHE[5][10] ), .C(\CACHE[6][10] ), 
        .D(\CACHE[7][10] ), .S0(n427), .S1(n441), .Y(n3121) );
  MXI4X1 U2204 ( .A(\CACHE[0][10] ), .B(\CACHE[1][10] ), .C(\CACHE[2][10] ), 
        .D(\CACHE[3][10] ), .S0(n427), .S1(n441), .Y(n3120) );
  MXI2X1 U2205 ( .A(n3122), .B(n3123), .S0(n464), .Y(N176) );
  MXI4X1 U2206 ( .A(\CACHE[4][11] ), .B(\CACHE[5][11] ), .C(\CACHE[6][11] ), 
        .D(\CACHE[7][11] ), .S0(n427), .S1(n441), .Y(n3123) );
  MXI4X1 U2207 ( .A(\CACHE[0][11] ), .B(\CACHE[1][11] ), .C(\CACHE[2][11] ), 
        .D(\CACHE[3][11] ), .S0(n427), .S1(n441), .Y(n3122) );
  MXI2X1 U2208 ( .A(n3124), .B(n3125), .S0(n465), .Y(N175) );
  MXI4X1 U2209 ( .A(\CACHE[4][12] ), .B(\CACHE[5][12] ), .C(\CACHE[6][12] ), 
        .D(\CACHE[7][12] ), .S0(n427), .S1(n442), .Y(n3125) );
  MXI4X1 U2210 ( .A(\CACHE[0][12] ), .B(\CACHE[1][12] ), .C(\CACHE[2][12] ), 
        .D(\CACHE[3][12] ), .S0(n427), .S1(n442), .Y(n3124) );
  MXI2X1 U2211 ( .A(n3126), .B(n3127), .S0(n465), .Y(N174) );
  MXI4X1 U2212 ( .A(\CACHE[4][13] ), .B(\CACHE[5][13] ), .C(\CACHE[6][13] ), 
        .D(\CACHE[7][13] ), .S0(n427), .S1(n442), .Y(n3127) );
  MXI4X1 U2213 ( .A(\CACHE[0][13] ), .B(\CACHE[1][13] ), .C(\CACHE[2][13] ), 
        .D(\CACHE[3][13] ), .S0(n427), .S1(n442), .Y(n3126) );
  MXI2X1 U2214 ( .A(n3128), .B(n3129), .S0(n465), .Y(N173) );
  MXI4X1 U2215 ( .A(\CACHE[4][14] ), .B(\CACHE[5][14] ), .C(\CACHE[6][14] ), 
        .D(\CACHE[7][14] ), .S0(n428), .S1(n442), .Y(n3129) );
  MXI4X1 U2216 ( .A(\CACHE[0][14] ), .B(\CACHE[1][14] ), .C(\CACHE[2][14] ), 
        .D(\CACHE[3][14] ), .S0(n428), .S1(n442), .Y(n3128) );
  MXI2X1 U2217 ( .A(n3130), .B(n3131), .S0(n465), .Y(N172) );
  MXI4X1 U2218 ( .A(\CACHE[4][15] ), .B(\CACHE[5][15] ), .C(\CACHE[6][15] ), 
        .D(\CACHE[7][15] ), .S0(n428), .S1(n442), .Y(n3131) );
  MXI4X1 U2219 ( .A(\CACHE[0][15] ), .B(\CACHE[1][15] ), .C(\CACHE[2][15] ), 
        .D(\CACHE[3][15] ), .S0(n428), .S1(n442), .Y(n3130) );
  MXI2X1 U2220 ( .A(n3132), .B(n3133), .S0(n465), .Y(N171) );
  MXI4X1 U2221 ( .A(\CACHE[4][16] ), .B(\CACHE[5][16] ), .C(\CACHE[6][16] ), 
        .D(\CACHE[7][16] ), .S0(n428), .S1(n442), .Y(n3133) );
  MXI4X1 U2222 ( .A(\CACHE[0][16] ), .B(\CACHE[1][16] ), .C(\CACHE[2][16] ), 
        .D(\CACHE[3][16] ), .S0(n428), .S1(n442), .Y(n3132) );
  MXI2X1 U2223 ( .A(n3134), .B(n3135), .S0(n465), .Y(N170) );
  MXI4X1 U2224 ( .A(\CACHE[4][17] ), .B(\CACHE[5][17] ), .C(\CACHE[6][17] ), 
        .D(\CACHE[7][17] ), .S0(n428), .S1(n442), .Y(n3135) );
  MXI4X1 U2225 ( .A(\CACHE[0][17] ), .B(\CACHE[1][17] ), .C(\CACHE[2][17] ), 
        .D(\CACHE[3][17] ), .S0(n428), .S1(n442), .Y(n3134) );
  MXI2X1 U2226 ( .A(n3136), .B(n3137), .S0(n465), .Y(N169) );
  MXI4X1 U2227 ( .A(\CACHE[4][18] ), .B(\CACHE[5][18] ), .C(\CACHE[6][18] ), 
        .D(\CACHE[7][18] ), .S0(n428), .S1(n443), .Y(n3137) );
  MXI4X1 U2228 ( .A(\CACHE[0][18] ), .B(\CACHE[1][18] ), .C(\CACHE[2][18] ), 
        .D(\CACHE[3][18] ), .S0(n428), .S1(n443), .Y(n3136) );
  MXI2X1 U2229 ( .A(n3138), .B(n3139), .S0(n465), .Y(N168) );
  MXI4X1 U2230 ( .A(\CACHE[4][19] ), .B(\CACHE[5][19] ), .C(\CACHE[6][19] ), 
        .D(\CACHE[7][19] ), .S0(n428), .S1(n443), .Y(n3139) );
  MXI4X1 U2231 ( .A(\CACHE[0][19] ), .B(\CACHE[1][19] ), .C(\CACHE[2][19] ), 
        .D(\CACHE[3][19] ), .S0(n428), .S1(n443), .Y(n3138) );
  MXI2X1 U2232 ( .A(n3140), .B(n3141), .S0(n465), .Y(N167) );
  MXI4X1 U2233 ( .A(\CACHE[4][20] ), .B(\CACHE[5][20] ), .C(\CACHE[6][20] ), 
        .D(\CACHE[7][20] ), .S0(n428), .S1(n443), .Y(n3141) );
  MXI4X1 U2234 ( .A(\CACHE[0][20] ), .B(\CACHE[1][20] ), .C(\CACHE[2][20] ), 
        .D(\CACHE[3][20] ), .S0(n429), .S1(n443), .Y(n3140) );
  MXI2X1 U2235 ( .A(n3142), .B(n3143), .S0(n465), .Y(N166) );
  MXI4X1 U2236 ( .A(\CACHE[4][21] ), .B(\CACHE[5][21] ), .C(\CACHE[6][21] ), 
        .D(\CACHE[7][21] ), .S0(n429), .S1(n443), .Y(n3143) );
  MXI4X1 U2237 ( .A(\CACHE[0][21] ), .B(\CACHE[1][21] ), .C(\CACHE[2][21] ), 
        .D(\CACHE[3][21] ), .S0(n429), .S1(n443), .Y(n3142) );
  MXI2X1 U2238 ( .A(n3144), .B(n3145), .S0(n465), .Y(N165) );
  MXI4X1 U2239 ( .A(\CACHE[4][22] ), .B(\CACHE[5][22] ), .C(\CACHE[6][22] ), 
        .D(\CACHE[7][22] ), .S0(n429), .S1(n443), .Y(n3145) );
  MXI4X1 U2240 ( .A(\CACHE[0][22] ), .B(\CACHE[1][22] ), .C(\CACHE[2][22] ), 
        .D(\CACHE[3][22] ), .S0(n429), .S1(n443), .Y(n3144) );
  MXI2X1 U2241 ( .A(n3146), .B(n3147), .S0(n465), .Y(N164) );
  MXI4X1 U2242 ( .A(\CACHE[4][23] ), .B(\CACHE[5][23] ), .C(\CACHE[6][23] ), 
        .D(\CACHE[7][23] ), .S0(n429), .S1(n443), .Y(n3147) );
  MXI4X1 U2243 ( .A(\CACHE[0][23] ), .B(\CACHE[1][23] ), .C(\CACHE[2][23] ), 
        .D(\CACHE[3][23] ), .S0(n429), .S1(n443), .Y(n3146) );
  MXI2X1 U2244 ( .A(n3148), .B(n3149), .S0(n466), .Y(N163) );
  MXI4X1 U2245 ( .A(\CACHE[4][24] ), .B(\CACHE[5][24] ), .C(\CACHE[6][24] ), 
        .D(\CACHE[7][24] ), .S0(n429), .S1(n444), .Y(n3149) );
  MXI4X1 U2246 ( .A(\CACHE[0][24] ), .B(\CACHE[1][24] ), .C(\CACHE[2][24] ), 
        .D(\CACHE[3][24] ), .S0(n429), .S1(n444), .Y(n3148) );
  MXI2X1 U2247 ( .A(n3150), .B(n3151), .S0(n466), .Y(N162) );
  MXI4X1 U2248 ( .A(\CACHE[4][25] ), .B(\CACHE[5][25] ), .C(\CACHE[6][25] ), 
        .D(\CACHE[7][25] ), .S0(n429), .S1(n444), .Y(n3151) );
  MXI4X1 U2249 ( .A(\CACHE[0][25] ), .B(\CACHE[1][25] ), .C(\CACHE[2][25] ), 
        .D(\CACHE[3][25] ), .S0(n429), .S1(n444), .Y(n3150) );
  MXI2X1 U2250 ( .A(n3152), .B(n3153), .S0(n466), .Y(N161) );
  MXI4X1 U2251 ( .A(\CACHE[4][26] ), .B(\CACHE[5][26] ), .C(\CACHE[6][26] ), 
        .D(\CACHE[7][26] ), .S0(n429), .S1(n444), .Y(n3153) );
  MXI4X1 U2252 ( .A(\CACHE[0][26] ), .B(\CACHE[1][26] ), .C(\CACHE[2][26] ), 
        .D(\CACHE[3][26] ), .S0(n429), .S1(n444), .Y(n3152) );
  MXI2X1 U2253 ( .A(n3154), .B(n3155), .S0(n466), .Y(N160) );
  MXI4X1 U2254 ( .A(\CACHE[4][27] ), .B(\CACHE[5][27] ), .C(\CACHE[6][27] ), 
        .D(\CACHE[7][27] ), .S0(n424), .S1(n444), .Y(n3155) );
  MXI4X1 U2255 ( .A(\CACHE[0][27] ), .B(\CACHE[1][27] ), .C(\CACHE[2][27] ), 
        .D(\CACHE[3][27] ), .S0(n429), .S1(n444), .Y(n3154) );
  MXI2X1 U2256 ( .A(n3156), .B(n3157), .S0(n466), .Y(N159) );
  MXI4X1 U2257 ( .A(\CACHE[4][28] ), .B(\CACHE[5][28] ), .C(\CACHE[6][28] ), 
        .D(\CACHE[7][28] ), .S0(N30), .S1(n444), .Y(n3157) );
  MXI4X1 U2258 ( .A(\CACHE[0][28] ), .B(\CACHE[1][28] ), .C(\CACHE[2][28] ), 
        .D(\CACHE[3][28] ), .S0(n425), .S1(n444), .Y(n3156) );
  MXI2X1 U2259 ( .A(n3158), .B(n3159), .S0(n466), .Y(N158) );
  MXI4X1 U2260 ( .A(\CACHE[4][29] ), .B(\CACHE[5][29] ), .C(\CACHE[6][29] ), 
        .D(\CACHE[7][29] ), .S0(N30), .S1(n444), .Y(n3159) );
  MXI4X1 U2261 ( .A(\CACHE[0][29] ), .B(\CACHE[1][29] ), .C(\CACHE[2][29] ), 
        .D(\CACHE[3][29] ), .S0(N30), .S1(n444), .Y(n3158) );
  MXI2X1 U2262 ( .A(n3160), .B(n3161), .S0(n466), .Y(N157) );
  MXI4X1 U2263 ( .A(\CACHE[4][30] ), .B(\CACHE[5][30] ), .C(\CACHE[6][30] ), 
        .D(\CACHE[7][30] ), .S0(N30), .S1(n440), .Y(n3161) );
  MXI4X1 U2264 ( .A(\CACHE[0][30] ), .B(\CACHE[1][30] ), .C(\CACHE[2][30] ), 
        .D(\CACHE[3][30] ), .S0(N30), .S1(n445), .Y(n3160) );
  MXI2X1 U2265 ( .A(n3162), .B(n3163), .S0(n466), .Y(N156) );
  MXI4X1 U2266 ( .A(\CACHE[4][31] ), .B(\CACHE[5][31] ), .C(\CACHE[6][31] ), 
        .D(\CACHE[7][31] ), .S0(N30), .S1(n456), .Y(n3163) );
  MXI4X1 U2267 ( .A(\CACHE[0][31] ), .B(\CACHE[1][31] ), .C(\CACHE[2][31] ), 
        .D(\CACHE[3][31] ), .S0(N30), .S1(n442), .Y(n3162) );
  MXI2X1 U2268 ( .A(n3164), .B(n3165), .S0(n466), .Y(N155) );
  MXI4X1 U2269 ( .A(\CACHE[4][32] ), .B(\CACHE[5][32] ), .C(\CACHE[6][32] ), 
        .D(\CACHE[7][32] ), .S0(N30), .S1(n447), .Y(n3165) );
  MXI4X1 U2270 ( .A(\CACHE[0][32] ), .B(\CACHE[1][32] ), .C(\CACHE[2][32] ), 
        .D(\CACHE[3][32] ), .S0(N30), .S1(n452), .Y(n3164) );
  MXI2X1 U2271 ( .A(n3166), .B(n3167), .S0(n466), .Y(N154) );
  MXI4X1 U2272 ( .A(\CACHE[4][33] ), .B(\CACHE[5][33] ), .C(\CACHE[6][33] ), 
        .D(\CACHE[7][33] ), .S0(N30), .S1(n449), .Y(n3167) );
  MXI4X1 U2273 ( .A(\CACHE[0][33] ), .B(\CACHE[1][33] ), .C(\CACHE[2][33] ), 
        .D(\CACHE[3][33] ), .S0(n430), .S1(n448), .Y(n3166) );
  MXI2X1 U2274 ( .A(n3168), .B(n3169), .S0(n466), .Y(N153) );
  MXI4X1 U2275 ( .A(\CACHE[4][34] ), .B(\CACHE[5][34] ), .C(\CACHE[6][34] ), 
        .D(\CACHE[7][34] ), .S0(n430), .S1(n441), .Y(n3169) );
  MXI4X1 U2276 ( .A(\CACHE[0][34] ), .B(\CACHE[1][34] ), .C(\CACHE[2][34] ), 
        .D(\CACHE[3][34] ), .S0(n430), .S1(n458), .Y(n3168) );
  MXI2X1 U2277 ( .A(n3170), .B(n3171), .S0(n466), .Y(N152) );
  MXI4X1 U2278 ( .A(\CACHE[4][35] ), .B(\CACHE[5][35] ), .C(\CACHE[6][35] ), 
        .D(\CACHE[7][35] ), .S0(n430), .S1(n453), .Y(n3171) );
  MXI4X1 U2279 ( .A(\CACHE[0][35] ), .B(\CACHE[1][35] ), .C(\CACHE[2][35] ), 
        .D(\CACHE[3][35] ), .S0(n430), .S1(n454), .Y(n3170) );
  MXI2X1 U2280 ( .A(n3172), .B(n3173), .S0(n467), .Y(N151) );
  MXI4X1 U2281 ( .A(\CACHE[4][36] ), .B(\CACHE[5][36] ), .C(\CACHE[6][36] ), 
        .D(\CACHE[7][36] ), .S0(n430), .S1(n445), .Y(n3173) );
  MXI4X1 U2282 ( .A(\CACHE[0][36] ), .B(\CACHE[1][36] ), .C(\CACHE[2][36] ), 
        .D(\CACHE[3][36] ), .S0(n430), .S1(n445), .Y(n3172) );
  MXI2X1 U2283 ( .A(n3174), .B(n3175), .S0(n467), .Y(N150) );
  MXI4X1 U2284 ( .A(\CACHE[4][37] ), .B(\CACHE[5][37] ), .C(\CACHE[6][37] ), 
        .D(\CACHE[7][37] ), .S0(n430), .S1(n445), .Y(n3175) );
  MXI4X1 U2285 ( .A(\CACHE[0][37] ), .B(\CACHE[1][37] ), .C(\CACHE[2][37] ), 
        .D(\CACHE[3][37] ), .S0(n430), .S1(n445), .Y(n3174) );
  MXI2X1 U2286 ( .A(n3176), .B(n3177), .S0(n467), .Y(N149) );
  MXI4X1 U2287 ( .A(\CACHE[4][38] ), .B(\CACHE[5][38] ), .C(\CACHE[6][38] ), 
        .D(\CACHE[7][38] ), .S0(n430), .S1(n445), .Y(n3177) );
  MXI4X1 U2288 ( .A(\CACHE[0][38] ), .B(\CACHE[1][38] ), .C(\CACHE[2][38] ), 
        .D(\CACHE[3][38] ), .S0(n430), .S1(n445), .Y(n3176) );
  MXI2X1 U2289 ( .A(n3178), .B(n3179), .S0(n467), .Y(N148) );
  MXI4X1 U2290 ( .A(\CACHE[4][39] ), .B(\CACHE[5][39] ), .C(\CACHE[6][39] ), 
        .D(\CACHE[7][39] ), .S0(n430), .S1(n445), .Y(n3179) );
  MXI4X1 U2291 ( .A(\CACHE[0][39] ), .B(\CACHE[1][39] ), .C(\CACHE[2][39] ), 
        .D(\CACHE[3][39] ), .S0(n431), .S1(n445), .Y(n3178) );
  MXI2X1 U2292 ( .A(n3180), .B(n3181), .S0(n467), .Y(N147) );
  MXI4X1 U2293 ( .A(\CACHE[4][40] ), .B(\CACHE[5][40] ), .C(\CACHE[6][40] ), 
        .D(\CACHE[7][40] ), .S0(n431), .S1(n445), .Y(n3181) );
  MXI4X1 U2294 ( .A(\CACHE[0][40] ), .B(\CACHE[1][40] ), .C(\CACHE[2][40] ), 
        .D(\CACHE[3][40] ), .S0(n431), .S1(n445), .Y(n3180) );
  MXI2X1 U2295 ( .A(n3182), .B(n3183), .S0(n467), .Y(N146) );
  MXI4X1 U2296 ( .A(\CACHE[4][41] ), .B(\CACHE[5][41] ), .C(\CACHE[6][41] ), 
        .D(\CACHE[7][41] ), .S0(n431), .S1(n445), .Y(n3183) );
  MXI4X1 U2297 ( .A(\CACHE[0][41] ), .B(\CACHE[1][41] ), .C(\CACHE[2][41] ), 
        .D(\CACHE[3][41] ), .S0(n431), .S1(n445), .Y(n3182) );
  MXI2X1 U2298 ( .A(n3184), .B(n3185), .S0(n467), .Y(N145) );
  MXI4X1 U2299 ( .A(\CACHE[4][42] ), .B(\CACHE[5][42] ), .C(\CACHE[6][42] ), 
        .D(\CACHE[7][42] ), .S0(n431), .S1(n453), .Y(n3185) );
  MXI4X1 U2300 ( .A(\CACHE[0][42] ), .B(\CACHE[1][42] ), .C(\CACHE[2][42] ), 
        .D(\CACHE[3][42] ), .S0(n431), .S1(n454), .Y(n3184) );
  MXI2X1 U2301 ( .A(n3186), .B(n3187), .S0(n467), .Y(N144) );
  MXI4X1 U2302 ( .A(\CACHE[4][43] ), .B(\CACHE[5][43] ), .C(\CACHE[6][43] ), 
        .D(\CACHE[7][43] ), .S0(n431), .S1(n450), .Y(n3187) );
  MXI4X1 U2303 ( .A(\CACHE[0][43] ), .B(\CACHE[1][43] ), .C(\CACHE[2][43] ), 
        .D(\CACHE[3][43] ), .S0(n431), .S1(n445), .Y(n3186) );
  MXI2X1 U2304 ( .A(n3188), .B(n3189), .S0(n467), .Y(N143) );
  MXI4X1 U2305 ( .A(\CACHE[4][44] ), .B(\CACHE[5][44] ), .C(\CACHE[6][44] ), 
        .D(\CACHE[7][44] ), .S0(n431), .S1(n446), .Y(n3189) );
  MXI4X1 U2306 ( .A(\CACHE[0][44] ), .B(\CACHE[1][44] ), .C(\CACHE[2][44] ), 
        .D(\CACHE[3][44] ), .S0(n431), .S1(n451), .Y(n3188) );
  MXI2X1 U2307 ( .A(n3190), .B(n3191), .S0(n467), .Y(N142) );
  MXI4X1 U2308 ( .A(\CACHE[4][45] ), .B(\CACHE[5][45] ), .C(\CACHE[6][45] ), 
        .D(\CACHE[7][45] ), .S0(n431), .S1(n457), .Y(n3191) );
  MXI4X1 U2309 ( .A(\CACHE[0][45] ), .B(\CACHE[1][45] ), .C(\CACHE[2][45] ), 
        .D(\CACHE[3][45] ), .S0(n431), .S1(n455), .Y(n3190) );
  MXI2X1 U2310 ( .A(n3192), .B(n3193), .S0(n467), .Y(N141) );
  MXI4X1 U2311 ( .A(\CACHE[4][46] ), .B(\CACHE[5][46] ), .C(\CACHE[6][46] ), 
        .D(\CACHE[7][46] ), .S0(n432), .S1(n459), .Y(n3193) );
  MXI4X1 U2312 ( .A(\CACHE[0][46] ), .B(\CACHE[1][46] ), .C(\CACHE[2][46] ), 
        .D(\CACHE[3][46] ), .S0(n432), .S1(n456), .Y(n3192) );
  MXI2X1 U2313 ( .A(n3194), .B(n3195), .S0(n467), .Y(N140) );
  MXI4X1 U2314 ( .A(\CACHE[4][47] ), .B(\CACHE[5][47] ), .C(\CACHE[6][47] ), 
        .D(\CACHE[7][47] ), .S0(n432), .S1(n444), .Y(n3195) );
  MXI4X1 U2315 ( .A(\CACHE[0][47] ), .B(\CACHE[1][47] ), .C(\CACHE[2][47] ), 
        .D(\CACHE[3][47] ), .S0(n432), .S1(n443), .Y(n3194) );
  MXI2X1 U2316 ( .A(n3196), .B(n3197), .S0(n468), .Y(N139) );
  MXI4X1 U2317 ( .A(\CACHE[4][48] ), .B(\CACHE[5][48] ), .C(\CACHE[6][48] ), 
        .D(\CACHE[7][48] ), .S0(n432), .S1(n446), .Y(n3197) );
  MXI4X1 U2318 ( .A(\CACHE[0][48] ), .B(\CACHE[1][48] ), .C(\CACHE[2][48] ), 
        .D(\CACHE[3][48] ), .S0(n432), .S1(n446), .Y(n3196) );
  MXI2X1 U2319 ( .A(n3198), .B(n3199), .S0(n468), .Y(N138) );
  MXI4X1 U2320 ( .A(\CACHE[4][49] ), .B(\CACHE[5][49] ), .C(\CACHE[6][49] ), 
        .D(\CACHE[7][49] ), .S0(n432), .S1(n446), .Y(n3199) );
  MXI4X1 U2321 ( .A(\CACHE[0][49] ), .B(\CACHE[1][49] ), .C(\CACHE[2][49] ), 
        .D(\CACHE[3][49] ), .S0(n432), .S1(n446), .Y(n3198) );
  MXI2X1 U2322 ( .A(n3200), .B(n3201), .S0(n468), .Y(N137) );
  MXI4X1 U2323 ( .A(\CACHE[4][50] ), .B(\CACHE[5][50] ), .C(\CACHE[6][50] ), 
        .D(\CACHE[7][50] ), .S0(n432), .S1(n446), .Y(n3201) );
  MXI4X1 U2324 ( .A(\CACHE[0][50] ), .B(\CACHE[1][50] ), .C(\CACHE[2][50] ), 
        .D(\CACHE[3][50] ), .S0(n432), .S1(n446), .Y(n3200) );
  MXI2X1 U2325 ( .A(n3202), .B(n3203), .S0(n468), .Y(N136) );
  MXI4X1 U2326 ( .A(\CACHE[4][51] ), .B(\CACHE[5][51] ), .C(\CACHE[6][51] ), 
        .D(\CACHE[7][51] ), .S0(n432), .S1(n446), .Y(n3203) );
  MXI4X1 U2327 ( .A(\CACHE[0][51] ), .B(\CACHE[1][51] ), .C(\CACHE[2][51] ), 
        .D(\CACHE[3][51] ), .S0(n432), .S1(n446), .Y(n3202) );
  MXI2X1 U2328 ( .A(n3204), .B(n3205), .S0(n468), .Y(N135) );
  MXI4X1 U2329 ( .A(\CACHE[4][52] ), .B(\CACHE[5][52] ), .C(\CACHE[6][52] ), 
        .D(\CACHE[7][52] ), .S0(n433), .S1(n446), .Y(n3205) );
  MXI4X1 U2330 ( .A(\CACHE[0][52] ), .B(\CACHE[1][52] ), .C(\CACHE[2][52] ), 
        .D(\CACHE[3][52] ), .S0(n433), .S1(n446), .Y(n3204) );
  MXI2X1 U2331 ( .A(n3206), .B(n3207), .S0(n468), .Y(N134) );
  MXI4X1 U2332 ( .A(\CACHE[4][53] ), .B(\CACHE[5][53] ), .C(\CACHE[6][53] ), 
        .D(\CACHE[7][53] ), .S0(n432), .S1(n446), .Y(n3207) );
  MXI4X1 U2333 ( .A(\CACHE[0][53] ), .B(\CACHE[1][53] ), .C(\CACHE[2][53] ), 
        .D(\CACHE[3][53] ), .S0(n433), .S1(n446), .Y(n3206) );
  MXI2X1 U2334 ( .A(n3208), .B(n3209), .S0(n468), .Y(N133) );
  MXI4X1 U2335 ( .A(\CACHE[4][54] ), .B(\CACHE[5][54] ), .C(\CACHE[6][54] ), 
        .D(\CACHE[7][54] ), .S0(n433), .S1(n447), .Y(n3209) );
  MXI4X1 U2336 ( .A(\CACHE[0][54] ), .B(\CACHE[1][54] ), .C(\CACHE[2][54] ), 
        .D(\CACHE[3][54] ), .S0(n433), .S1(n447), .Y(n3208) );
  MXI2X1 U2337 ( .A(n3210), .B(n3211), .S0(n468), .Y(N132) );
  MXI4X1 U2338 ( .A(\CACHE[4][55] ), .B(\CACHE[5][55] ), .C(\CACHE[6][55] ), 
        .D(\CACHE[7][55] ), .S0(n433), .S1(n447), .Y(n3211) );
  MXI4X1 U2339 ( .A(\CACHE[0][55] ), .B(\CACHE[1][55] ), .C(\CACHE[2][55] ), 
        .D(\CACHE[3][55] ), .S0(n433), .S1(n447), .Y(n3210) );
  MXI2X1 U2340 ( .A(n3212), .B(n3213), .S0(n468), .Y(N131) );
  MXI4X1 U2341 ( .A(\CACHE[4][56] ), .B(\CACHE[5][56] ), .C(\CACHE[6][56] ), 
        .D(\CACHE[7][56] ), .S0(n433), .S1(n447), .Y(n3213) );
  MXI4X1 U2342 ( .A(\CACHE[0][56] ), .B(\CACHE[1][56] ), .C(\CACHE[2][56] ), 
        .D(\CACHE[3][56] ), .S0(n433), .S1(n447), .Y(n3212) );
  MXI2X1 U2343 ( .A(n3214), .B(n3215), .S0(n468), .Y(N130) );
  MXI4X1 U2344 ( .A(\CACHE[4][57] ), .B(\CACHE[5][57] ), .C(\CACHE[6][57] ), 
        .D(\CACHE[7][57] ), .S0(n433), .S1(n447), .Y(n3215) );
  MXI4X1 U2345 ( .A(\CACHE[0][57] ), .B(\CACHE[1][57] ), .C(\CACHE[2][57] ), 
        .D(\CACHE[3][57] ), .S0(n433), .S1(n447), .Y(n3214) );
  MXI2X1 U2346 ( .A(n3216), .B(n3217), .S0(n468), .Y(N129) );
  MXI4X1 U2347 ( .A(\CACHE[4][58] ), .B(\CACHE[5][58] ), .C(\CACHE[6][58] ), 
        .D(\CACHE[7][58] ), .S0(n433), .S1(n447), .Y(n3217) );
  MXI4X1 U2348 ( .A(\CACHE[0][58] ), .B(\CACHE[1][58] ), .C(\CACHE[2][58] ), 
        .D(\CACHE[3][58] ), .S0(n434), .S1(n447), .Y(n3216) );
  MXI2X1 U2349 ( .A(n3218), .B(n3219), .S0(n468), .Y(N128) );
  MXI4X1 U2350 ( .A(\CACHE[4][59] ), .B(\CACHE[5][59] ), .C(\CACHE[6][59] ), 
        .D(\CACHE[7][59] ), .S0(n433), .S1(n447), .Y(n3219) );
  MXI4X1 U2351 ( .A(\CACHE[0][59] ), .B(\CACHE[1][59] ), .C(\CACHE[2][59] ), 
        .D(\CACHE[3][59] ), .S0(n434), .S1(n447), .Y(n3218) );
  MXI2X1 U2352 ( .A(n3220), .B(n3221), .S0(n471), .Y(N127) );
  MXI4X1 U2353 ( .A(\CACHE[4][60] ), .B(\CACHE[5][60] ), .C(\CACHE[6][60] ), 
        .D(\CACHE[7][60] ), .S0(n434), .S1(n448), .Y(n3221) );
  MXI4X1 U2354 ( .A(\CACHE[0][60] ), .B(\CACHE[1][60] ), .C(\CACHE[2][60] ), 
        .D(\CACHE[3][60] ), .S0(n434), .S1(n448), .Y(n3220) );
  MXI2X1 U2355 ( .A(n3222), .B(n3223), .S0(n464), .Y(N126) );
  MXI4X1 U2356 ( .A(\CACHE[4][61] ), .B(\CACHE[5][61] ), .C(\CACHE[6][61] ), 
        .D(\CACHE[7][61] ), .S0(n434), .S1(n448), .Y(n3223) );
  MXI4X1 U2357 ( .A(\CACHE[0][61] ), .B(\CACHE[1][61] ), .C(\CACHE[2][61] ), 
        .D(\CACHE[3][61] ), .S0(n434), .S1(n448), .Y(n3222) );
  MXI2X1 U2358 ( .A(n3224), .B(n3225), .S0(n465), .Y(N125) );
  MXI4X1 U2359 ( .A(\CACHE[4][62] ), .B(\CACHE[5][62] ), .C(\CACHE[6][62] ), 
        .D(\CACHE[7][62] ), .S0(n434), .S1(n448), .Y(n3225) );
  MXI4X1 U2360 ( .A(\CACHE[0][62] ), .B(\CACHE[1][62] ), .C(\CACHE[2][62] ), 
        .D(\CACHE[3][62] ), .S0(n434), .S1(n448), .Y(n3224) );
  MXI2X1 U2361 ( .A(n3226), .B(n3227), .S0(n466), .Y(N124) );
  MXI4X1 U2362 ( .A(\CACHE[4][63] ), .B(\CACHE[5][63] ), .C(\CACHE[6][63] ), 
        .D(\CACHE[7][63] ), .S0(n434), .S1(n448), .Y(n3227) );
  MXI4X1 U2363 ( .A(\CACHE[0][63] ), .B(\CACHE[1][63] ), .C(\CACHE[2][63] ), 
        .D(\CACHE[3][63] ), .S0(n434), .S1(n448), .Y(n3226) );
  MXI2X1 U2364 ( .A(n3292), .B(n3293), .S0(n469), .Y(N91) );
  MXI4X1 U2365 ( .A(\CACHE[4][96] ), .B(\CACHE[5][96] ), .C(\CACHE[6][96] ), 
        .D(\CACHE[7][96] ), .S0(n433), .S1(n453), .Y(n3293) );
  MXI4X1 U2366 ( .A(\CACHE[0][96] ), .B(\CACHE[1][96] ), .C(\CACHE[2][96] ), 
        .D(\CACHE[3][96] ), .S0(n432), .S1(n453), .Y(n3292) );
  MXI2X1 U2367 ( .A(n3294), .B(n3295), .S0(n469), .Y(N90) );
  MXI4X1 U2368 ( .A(\CACHE[4][97] ), .B(\CACHE[5][97] ), .C(\CACHE[6][97] ), 
        .D(\CACHE[7][97] ), .S0(n422), .S1(n453), .Y(n3295) );
  MXI4X1 U2369 ( .A(\CACHE[0][97] ), .B(\CACHE[1][97] ), .C(\CACHE[2][97] ), 
        .D(\CACHE[3][97] ), .S0(n430), .S1(n453), .Y(n3294) );
  MXI2X1 U2370 ( .A(n3296), .B(n3297), .S0(n469), .Y(N89) );
  MXI4X1 U2371 ( .A(\CACHE[4][98] ), .B(\CACHE[5][98] ), .C(\CACHE[6][98] ), 
        .D(\CACHE[7][98] ), .S0(n428), .S1(n453), .Y(n3297) );
  MXI4X1 U2372 ( .A(\CACHE[0][98] ), .B(\CACHE[1][98] ), .C(\CACHE[2][98] ), 
        .D(\CACHE[3][98] ), .S0(n435), .S1(n453), .Y(n3296) );
  MXI2X1 U2373 ( .A(n3298), .B(n3299), .S0(n469), .Y(N88) );
  MXI4X1 U2374 ( .A(\CACHE[4][99] ), .B(\CACHE[5][99] ), .C(\CACHE[6][99] ), 
        .D(\CACHE[7][99] ), .S0(n434), .S1(n453), .Y(n3299) );
  MXI4X1 U2375 ( .A(\CACHE[0][99] ), .B(\CACHE[1][99] ), .C(\CACHE[2][99] ), 
        .D(\CACHE[3][99] ), .S0(n420), .S1(n453), .Y(n3298) );
  MXI2X1 U2376 ( .A(n3300), .B(n3301), .S0(n469), .Y(N87) );
  MXI4X1 U2377 ( .A(\CACHE[4][100] ), .B(\CACHE[5][100] ), .C(\CACHE[6][100] ), 
        .D(\CACHE[7][100] ), .S0(n418), .S1(n453), .Y(n3301) );
  MXI4X1 U2378 ( .A(\CACHE[0][100] ), .B(\CACHE[1][100] ), .C(\CACHE[2][100] ), 
        .D(\CACHE[3][100] ), .S0(n431), .S1(n453), .Y(n3300) );
  MXI2X1 U2379 ( .A(n3302), .B(n3303), .S0(n469), .Y(N86) );
  MXI4X1 U2380 ( .A(\CACHE[4][101] ), .B(\CACHE[5][101] ), .C(\CACHE[6][101] ), 
        .D(\CACHE[7][101] ), .S0(n426), .S1(n453), .Y(n3303) );
  MXI4X1 U2381 ( .A(\CACHE[0][101] ), .B(\CACHE[1][101] ), .C(\CACHE[2][101] ), 
        .D(\CACHE[3][101] ), .S0(n419), .S1(n453), .Y(n3302) );
  MXI2X1 U2382 ( .A(n3304), .B(n3305), .S0(n469), .Y(N85) );
  MXI4X1 U2383 ( .A(\CACHE[4][102] ), .B(\CACHE[5][102] ), .C(\CACHE[6][102] ), 
        .D(\CACHE[7][102] ), .S0(n424), .S1(n454), .Y(n3305) );
  MXI4X1 U2384 ( .A(\CACHE[0][102] ), .B(\CACHE[1][102] ), .C(\CACHE[2][102] ), 
        .D(\CACHE[3][102] ), .S0(n429), .S1(n454), .Y(n3304) );
  MXI2X1 U2385 ( .A(n3306), .B(n3307), .S0(n469), .Y(N84) );
  MXI4X1 U2386 ( .A(\CACHE[4][103] ), .B(\CACHE[5][103] ), .C(\CACHE[6][103] ), 
        .D(\CACHE[7][103] ), .S0(n425), .S1(n454), .Y(n3307) );
  MXI4X1 U2387 ( .A(\CACHE[0][103] ), .B(\CACHE[1][103] ), .C(\CACHE[2][103] ), 
        .D(\CACHE[3][103] ), .S0(n420), .S1(n454), .Y(n3306) );
  MXI2X1 U2388 ( .A(n3308), .B(n3309), .S0(n469), .Y(N83) );
  MXI4X1 U2389 ( .A(\CACHE[4][104] ), .B(\CACHE[5][104] ), .C(\CACHE[6][104] ), 
        .D(\CACHE[7][104] ), .S0(n420), .S1(n454), .Y(n3309) );
  MXI4X1 U2390 ( .A(\CACHE[0][104] ), .B(\CACHE[1][104] ), .C(\CACHE[2][104] ), 
        .D(\CACHE[3][104] ), .S0(n420), .S1(n454), .Y(n3308) );
  MXI2X1 U2391 ( .A(n3310), .B(n3311), .S0(n469), .Y(N82) );
  MXI4X1 U2392 ( .A(\CACHE[4][105] ), .B(\CACHE[5][105] ), .C(\CACHE[6][105] ), 
        .D(\CACHE[7][105] ), .S0(n420), .S1(n454), .Y(n3311) );
  MXI4X1 U2393 ( .A(\CACHE[0][105] ), .B(\CACHE[1][105] ), .C(\CACHE[2][105] ), 
        .D(\CACHE[3][105] ), .S0(n420), .S1(n454), .Y(n3310) );
  MXI2X1 U2394 ( .A(n3312), .B(n3313), .S0(n469), .Y(N81) );
  MXI4X1 U2395 ( .A(\CACHE[4][106] ), .B(\CACHE[5][106] ), .C(\CACHE[6][106] ), 
        .D(\CACHE[7][106] ), .S0(n420), .S1(n454), .Y(n3313) );
  MXI4X1 U2396 ( .A(\CACHE[0][106] ), .B(\CACHE[1][106] ), .C(\CACHE[2][106] ), 
        .D(\CACHE[3][106] ), .S0(n420), .S1(n454), .Y(n3312) );
  MXI2X1 U2397 ( .A(n3314), .B(n3315), .S0(n469), .Y(N80) );
  MXI4X1 U2398 ( .A(\CACHE[4][107] ), .B(\CACHE[5][107] ), .C(\CACHE[6][107] ), 
        .D(\CACHE[7][107] ), .S0(n420), .S1(n454), .Y(n3315) );
  MXI4X1 U2399 ( .A(\CACHE[0][107] ), .B(\CACHE[1][107] ), .C(\CACHE[2][107] ), 
        .D(\CACHE[3][107] ), .S0(n420), .S1(n454), .Y(n3314) );
  MXI2X1 U2400 ( .A(n3316), .B(n3317), .S0(n470), .Y(N79) );
  MXI4X1 U2401 ( .A(\CACHE[4][108] ), .B(\CACHE[5][108] ), .C(\CACHE[6][108] ), 
        .D(\CACHE[7][108] ), .S0(n420), .S1(n455), .Y(n3317) );
  MXI4X1 U2402 ( .A(\CACHE[0][108] ), .B(\CACHE[1][108] ), .C(\CACHE[2][108] ), 
        .D(\CACHE[3][108] ), .S0(n420), .S1(n455), .Y(n3316) );
  MXI2X1 U2403 ( .A(n3318), .B(n3319), .S0(n470), .Y(N78) );
  MXI4X1 U2404 ( .A(\CACHE[4][109] ), .B(\CACHE[5][109] ), .C(\CACHE[6][109] ), 
        .D(\CACHE[7][109] ), .S0(n420), .S1(n455), .Y(n3319) );
  MXI4X1 U2405 ( .A(\CACHE[0][109] ), .B(\CACHE[1][109] ), .C(\CACHE[2][109] ), 
        .D(\CACHE[3][109] ), .S0(n420), .S1(n455), .Y(n3318) );
  MXI2X1 U2406 ( .A(n3320), .B(n3321), .S0(n470), .Y(N77) );
  MXI4X1 U2407 ( .A(\CACHE[4][110] ), .B(\CACHE[5][110] ), .C(\CACHE[6][110] ), 
        .D(\CACHE[7][110] ), .S0(n422), .S1(n455), .Y(n3321) );
  MXI4X1 U2408 ( .A(\CACHE[0][110] ), .B(\CACHE[1][110] ), .C(\CACHE[2][110] ), 
        .D(\CACHE[3][110] ), .S0(n430), .S1(n455), .Y(n3320) );
  MXI2X1 U2409 ( .A(n3322), .B(n3323), .S0(n470), .Y(N76) );
  MXI4X1 U2410 ( .A(\CACHE[4][111] ), .B(\CACHE[5][111] ), .C(\CACHE[6][111] ), 
        .D(\CACHE[7][111] ), .S0(n434), .S1(n455), .Y(n3323) );
  MXI4X1 U2411 ( .A(\CACHE[0][111] ), .B(\CACHE[1][111] ), .C(\CACHE[2][111] ), 
        .D(\CACHE[3][111] ), .S0(n420), .S1(n455), .Y(n3322) );
  MXI2X1 U2412 ( .A(n3324), .B(n3325), .S0(n470), .Y(N75) );
  MXI4X1 U2413 ( .A(\CACHE[4][112] ), .B(\CACHE[5][112] ), .C(\CACHE[6][112] ), 
        .D(\CACHE[7][112] ), .S0(n418), .S1(n455), .Y(n3325) );
  MXI4X1 U2414 ( .A(\CACHE[0][112] ), .B(\CACHE[1][112] ), .C(\CACHE[2][112] ), 
        .D(\CACHE[3][112] ), .S0(n431), .S1(n455), .Y(n3324) );
  MXI2X1 U2415 ( .A(n3326), .B(n3327), .S0(n470), .Y(N74) );
  MXI4X1 U2416 ( .A(\CACHE[4][113] ), .B(\CACHE[5][113] ), .C(\CACHE[6][113] ), 
        .D(\CACHE[7][113] ), .S0(n426), .S1(n455), .Y(n3327) );
  MXI4X1 U2417 ( .A(\CACHE[0][113] ), .B(\CACHE[1][113] ), .C(\CACHE[2][113] ), 
        .D(\CACHE[3][113] ), .S0(n419), .S1(n455), .Y(n3326) );
  MXI2X1 U2418 ( .A(n3328), .B(n3329), .S0(n470), .Y(N73) );
  MXI4X1 U2419 ( .A(\CACHE[4][114] ), .B(\CACHE[5][114] ), .C(\CACHE[6][114] ), 
        .D(\CACHE[7][114] ), .S0(n423), .S1(n456), .Y(n3329) );
  MXI4X1 U2420 ( .A(\CACHE[0][114] ), .B(\CACHE[1][114] ), .C(\CACHE[2][114] ), 
        .D(\CACHE[3][114] ), .S0(n421), .S1(n456), .Y(n3328) );
  MXI2X1 U2421 ( .A(n3330), .B(n3331), .S0(n470), .Y(N72) );
  MXI4X1 U2422 ( .A(\CACHE[4][115] ), .B(\CACHE[5][115] ), .C(\CACHE[6][115] ), 
        .D(\CACHE[7][115] ), .S0(n423), .S1(n456), .Y(n3331) );
  MXI4X1 U2423 ( .A(\CACHE[0][115] ), .B(\CACHE[1][115] ), .C(\CACHE[2][115] ), 
        .D(\CACHE[3][115] ), .S0(n427), .S1(n456), .Y(n3330) );
  MXI2X1 U2424 ( .A(n3332), .B(n3333), .S0(n470), .Y(N71) );
  MXI4X1 U2425 ( .A(\CACHE[4][116] ), .B(\CACHE[5][116] ), .C(\CACHE[6][116] ), 
        .D(\CACHE[7][116] ), .S0(n421), .S1(n456), .Y(n3333) );
  MXI4X1 U2426 ( .A(\CACHE[0][116] ), .B(\CACHE[1][116] ), .C(\CACHE[2][116] ), 
        .D(\CACHE[3][116] ), .S0(n421), .S1(n456), .Y(n3332) );
  MXI2X1 U2427 ( .A(n3334), .B(n3335), .S0(n470), .Y(N70) );
  MXI4X1 U2428 ( .A(\CACHE[4][117] ), .B(\CACHE[5][117] ), .C(\CACHE[6][117] ), 
        .D(\CACHE[7][117] ), .S0(n421), .S1(n456), .Y(n3335) );
  MXI4X1 U2429 ( .A(\CACHE[0][117] ), .B(\CACHE[1][117] ), .C(\CACHE[2][117] ), 
        .D(\CACHE[3][117] ), .S0(n418), .S1(n456), .Y(n3334) );
  MXI2X1 U2430 ( .A(n3336), .B(n3337), .S0(n470), .Y(N69) );
  MXI4X1 U2431 ( .A(\CACHE[4][118] ), .B(\CACHE[5][118] ), .C(\CACHE[6][118] ), 
        .D(\CACHE[7][118] ), .S0(n421), .S1(n456), .Y(n3337) );
  MXI4X1 U2432 ( .A(\CACHE[0][118] ), .B(\CACHE[1][118] ), .C(\CACHE[2][118] ), 
        .D(\CACHE[3][118] ), .S0(n421), .S1(n456), .Y(n3336) );
  MXI2X1 U2433 ( .A(n3338), .B(n3339), .S0(n470), .Y(N68) );
  MXI4X1 U2434 ( .A(\CACHE[4][119] ), .B(\CACHE[5][119] ), .C(\CACHE[6][119] ), 
        .D(\CACHE[7][119] ), .S0(n421), .S1(n456), .Y(n3339) );
  MXI4X1 U2435 ( .A(\CACHE[0][119] ), .B(\CACHE[1][119] ), .C(\CACHE[2][119] ), 
        .D(\CACHE[3][119] ), .S0(n421), .S1(n456), .Y(n3338) );
  MXI2X1 U2436 ( .A(n3340), .B(n3341), .S0(n471), .Y(N67) );
  MXI4X1 U2437 ( .A(\CACHE[4][120] ), .B(\CACHE[5][120] ), .C(\CACHE[6][120] ), 
        .D(\CACHE[7][120] ), .S0(n421), .S1(n452), .Y(n3341) );
  MXI4X1 U2438 ( .A(\CACHE[0][120] ), .B(\CACHE[1][120] ), .C(\CACHE[2][120] ), 
        .D(\CACHE[3][120] ), .S0(n421), .S1(n456), .Y(n3340) );
  MXI2X1 U2439 ( .A(n3342), .B(n3343), .S0(n467), .Y(N66) );
  MXI4X1 U2440 ( .A(\CACHE[4][121] ), .B(\CACHE[5][121] ), .C(\CACHE[6][121] ), 
        .D(\CACHE[7][121] ), .S0(n421), .S1(n448), .Y(n3343) );
  MXI4X1 U2441 ( .A(\CACHE[0][121] ), .B(\CACHE[1][121] ), .C(\CACHE[2][121] ), 
        .D(\CACHE[3][121] ), .S0(n421), .S1(n447), .Y(n3342) );
  MXI2X1 U2442 ( .A(n3344), .B(n3345), .S0(n468), .Y(N65) );
  MXI4X1 U2443 ( .A(\CACHE[4][122] ), .B(\CACHE[5][122] ), .C(\CACHE[6][122] ), 
        .D(\CACHE[7][122] ), .S0(n421), .S1(n460), .Y(n3345) );
  MXI4X1 U2444 ( .A(\CACHE[0][122] ), .B(\CACHE[1][122] ), .C(\CACHE[2][122] ), 
        .D(\CACHE[3][122] ), .S0(n421), .S1(n449), .Y(n3344) );
  MXI2X1 U2445 ( .A(n3346), .B(n3347), .S0(n464), .Y(N64) );
  MXI4X1 U2446 ( .A(\CACHE[4][123] ), .B(\CACHE[5][123] ), .C(\CACHE[6][123] ), 
        .D(\CACHE[7][123] ), .S0(n422), .S1(n453), .Y(n3347) );
  MXI4X1 U2447 ( .A(\CACHE[0][123] ), .B(\CACHE[1][123] ), .C(\CACHE[2][123] ), 
        .D(\CACHE[3][123] ), .S0(n422), .S1(n454), .Y(n3346) );
  MXI2X1 U2448 ( .A(n3348), .B(n3349), .S0(n465), .Y(N63) );
  MXI4X1 U2449 ( .A(\CACHE[4][124] ), .B(\CACHE[5][124] ), .C(\CACHE[6][124] ), 
        .D(\CACHE[7][124] ), .S0(n422), .S1(n440), .Y(n3349) );
  MXI4X1 U2450 ( .A(\CACHE[0][124] ), .B(\CACHE[1][124] ), .C(\CACHE[2][124] ), 
        .D(\CACHE[3][124] ), .S0(n422), .S1(n445), .Y(n3348) );
  MXI2X1 U2451 ( .A(n3350), .B(n3351), .S0(n466), .Y(N62) );
  MXI4X1 U2452 ( .A(\CACHE[4][125] ), .B(\CACHE[5][125] ), .C(\CACHE[6][125] ), 
        .D(\CACHE[7][125] ), .S0(n422), .S1(n450), .Y(n3351) );
  MXI4X1 U2453 ( .A(\CACHE[0][125] ), .B(\CACHE[1][125] ), .C(\CACHE[2][125] ), 
        .D(\CACHE[3][125] ), .S0(n422), .S1(n442), .Y(n3350) );
  MXI2X1 U2454 ( .A(n3352), .B(n3353), .S0(n469), .Y(N61) );
  MXI4X1 U2455 ( .A(\CACHE[4][126] ), .B(\CACHE[5][126] ), .C(\CACHE[6][126] ), 
        .D(\CACHE[7][126] ), .S0(n422), .S1(n457), .Y(n3353) );
  MXI4X1 U2456 ( .A(\CACHE[0][126] ), .B(\CACHE[1][126] ), .C(\CACHE[2][126] ), 
        .D(\CACHE[3][126] ), .S0(n422), .S1(n457), .Y(n3352) );
  MXI2X1 U2457 ( .A(n3354), .B(n3355), .S0(n470), .Y(N60) );
  MXI4X1 U2458 ( .A(\CACHE[4][127] ), .B(\CACHE[5][127] ), .C(\CACHE[6][127] ), 
        .D(\CACHE[7][127] ), .S0(n422), .S1(n457), .Y(n3355) );
  MXI4X1 U2459 ( .A(\CACHE[0][127] ), .B(\CACHE[1][127] ), .C(\CACHE[2][127] ), 
        .D(\CACHE[3][127] ), .S0(n422), .S1(n457), .Y(n3354) );
  MXI2X1 U2460 ( .A(n3228), .B(n3229), .S0(n469), .Y(N123) );
  MXI4X1 U2461 ( .A(\CACHE[4][64] ), .B(\CACHE[5][64] ), .C(\CACHE[6][64] ), 
        .D(\CACHE[7][64] ), .S0(n434), .S1(n448), .Y(n3229) );
  MXI4X1 U2462 ( .A(\CACHE[0][64] ), .B(\CACHE[1][64] ), .C(\CACHE[2][64] ), 
        .D(\CACHE[3][64] ), .S0(n434), .S1(n448), .Y(n3228) );
  MXI2X1 U2463 ( .A(n3230), .B(n3231), .S0(n470), .Y(N122) );
  MXI4X1 U2464 ( .A(\CACHE[4][65] ), .B(\CACHE[5][65] ), .C(\CACHE[6][65] ), 
        .D(\CACHE[7][65] ), .S0(n434), .S1(n448), .Y(n3231) );
  MXI4X1 U2465 ( .A(\CACHE[0][65] ), .B(\CACHE[1][65] ), .C(\CACHE[2][65] ), 
        .D(\CACHE[3][65] ), .S0(n435), .S1(n448), .Y(n3230) );
  MXI2X1 U2466 ( .A(n3232), .B(n3233), .S0(n467), .Y(N121) );
  MXI4X1 U2467 ( .A(\CACHE[4][66] ), .B(\CACHE[5][66] ), .C(\CACHE[6][66] ), 
        .D(\CACHE[7][66] ), .S0(n435), .S1(n449), .Y(n3233) );
  MXI4X1 U2468 ( .A(\CACHE[0][66] ), .B(\CACHE[1][66] ), .C(\CACHE[2][66] ), 
        .D(\CACHE[3][66] ), .S0(n435), .S1(n449), .Y(n3232) );
  MXI2X1 U2469 ( .A(n3234), .B(n3235), .S0(n467), .Y(N120) );
  MXI4X1 U2470 ( .A(\CACHE[4][67] ), .B(\CACHE[5][67] ), .C(\CACHE[6][67] ), 
        .D(\CACHE[7][67] ), .S0(n435), .S1(n449), .Y(n3235) );
  MXI4X1 U2471 ( .A(\CACHE[0][67] ), .B(\CACHE[1][67] ), .C(\CACHE[2][67] ), 
        .D(\CACHE[3][67] ), .S0(n435), .S1(n449), .Y(n3234) );
  MXI2X1 U2472 ( .A(n3236), .B(n3237), .S0(n468), .Y(N119) );
  MXI4X1 U2473 ( .A(\CACHE[4][68] ), .B(\CACHE[5][68] ), .C(\CACHE[6][68] ), 
        .D(\CACHE[7][68] ), .S0(n435), .S1(n449), .Y(n3237) );
  MXI4X1 U2474 ( .A(\CACHE[0][68] ), .B(\CACHE[1][68] ), .C(\CACHE[2][68] ), 
        .D(\CACHE[3][68] ), .S0(n435), .S1(n449), .Y(n3236) );
  MXI2X1 U2475 ( .A(n3238), .B(n3239), .S0(n472), .Y(N118) );
  MXI4X1 U2476 ( .A(\CACHE[4][69] ), .B(\CACHE[5][69] ), .C(\CACHE[6][69] ), 
        .D(\CACHE[7][69] ), .S0(n435), .S1(n449), .Y(n3239) );
  MXI4X1 U2477 ( .A(\CACHE[0][69] ), .B(\CACHE[1][69] ), .C(\CACHE[2][69] ), 
        .D(\CACHE[3][69] ), .S0(n435), .S1(n449), .Y(n3238) );
  MXI2X1 U2478 ( .A(n3240), .B(n3241), .S0(n471), .Y(N117) );
  MXI4X1 U2479 ( .A(\CACHE[4][70] ), .B(\CACHE[5][70] ), .C(\CACHE[6][70] ), 
        .D(\CACHE[7][70] ), .S0(n435), .S1(n449), .Y(n3241) );
  MXI4X1 U2480 ( .A(\CACHE[0][70] ), .B(\CACHE[1][70] ), .C(\CACHE[2][70] ), 
        .D(\CACHE[3][70] ), .S0(n435), .S1(n449), .Y(n3240) );
  MXI2X1 U2481 ( .A(n3242), .B(n3243), .S0(n464), .Y(N116) );
  MXI4X1 U2482 ( .A(\CACHE[4][71] ), .B(\CACHE[5][71] ), .C(\CACHE[6][71] ), 
        .D(\CACHE[7][71] ), .S0(n435), .S1(n449), .Y(n3243) );
  MXI4X1 U2483 ( .A(\CACHE[0][71] ), .B(\CACHE[1][71] ), .C(\CACHE[2][71] ), 
        .D(\CACHE[3][71] ), .S0(n436), .S1(n449), .Y(n3242) );
  MXI2X1 U2484 ( .A(n3244), .B(n3245), .S0(n468), .Y(N115) );
  MXI4X1 U2485 ( .A(\CACHE[4][72] ), .B(\CACHE[5][72] ), .C(\CACHE[6][72] ), 
        .D(\CACHE[7][72] ), .S0(n436), .S1(n447), .Y(n3245) );
  MXI4X1 U2486 ( .A(\CACHE[0][72] ), .B(\CACHE[1][72] ), .C(\CACHE[2][72] ), 
        .D(\CACHE[3][72] ), .S0(n435), .S1(n452), .Y(n3244) );
  MXI2X1 U2487 ( .A(n3246), .B(n3247), .S0(n472), .Y(N114) );
  MXI4X1 U2488 ( .A(\CACHE[4][73] ), .B(\CACHE[5][73] ), .C(\CACHE[6][73] ), 
        .D(\CACHE[7][73] ), .S0(n436), .S1(n449), .Y(n3247) );
  MXI4X1 U2489 ( .A(\CACHE[0][73] ), .B(\CACHE[1][73] ), .C(\CACHE[2][73] ), 
        .D(\CACHE[3][73] ), .S0(n436), .S1(n448), .Y(n3246) );
  MXI2X1 U2490 ( .A(n3248), .B(n3249), .S0(n472), .Y(N113) );
  MXI4X1 U2491 ( .A(\CACHE[4][74] ), .B(\CACHE[5][74] ), .C(\CACHE[6][74] ), 
        .D(\CACHE[7][74] ), .S0(n436), .S1(n441), .Y(n3249) );
  MXI4X1 U2492 ( .A(\CACHE[0][74] ), .B(\CACHE[1][74] ), .C(\CACHE[2][74] ), 
        .D(\CACHE[3][74] ), .S0(n436), .S1(n458), .Y(n3248) );
  MXI2X1 U2493 ( .A(n3250), .B(n3251), .S0(n471), .Y(N112) );
  MXI4X1 U2494 ( .A(\CACHE[4][75] ), .B(\CACHE[5][75] ), .C(\CACHE[6][75] ), 
        .D(\CACHE[7][75] ), .S0(n436), .S1(n455), .Y(n3251) );
  MXI4X1 U2495 ( .A(\CACHE[0][75] ), .B(\CACHE[1][75] ), .C(\CACHE[2][75] ), 
        .D(\CACHE[3][75] ), .S0(n436), .S1(n446), .Y(n3250) );
  MXI2X1 U2496 ( .A(n3252), .B(n3253), .S0(n464), .Y(N111) );
  MXI4X1 U2497 ( .A(\CACHE[4][76] ), .B(\CACHE[5][76] ), .C(\CACHE[6][76] ), 
        .D(\CACHE[7][76] ), .S0(n436), .S1(n459), .Y(n3253) );
  MXI4X1 U2498 ( .A(\CACHE[0][76] ), .B(\CACHE[1][76] ), .C(\CACHE[2][76] ), 
        .D(\CACHE[3][76] ), .S0(n436), .S1(n457), .Y(n3252) );
  MXI2X1 U2499 ( .A(n3254), .B(n3255), .S0(n465), .Y(N110) );
  MXI4X1 U2500 ( .A(\CACHE[4][77] ), .B(\CACHE[5][77] ), .C(\CACHE[6][77] ), 
        .D(\CACHE[7][77] ), .S0(n436), .S1(n444), .Y(n3255) );
  MXI4X1 U2501 ( .A(\CACHE[0][77] ), .B(\CACHE[1][77] ), .C(\CACHE[2][77] ), 
        .D(\CACHE[3][77] ), .S0(n436), .S1(n443), .Y(n3254) );
  MXI2X1 U2502 ( .A(n3256), .B(n3257), .S0(n466), .Y(N109) );
  MXI4X1 U2503 ( .A(\CACHE[4][78] ), .B(\CACHE[5][78] ), .C(\CACHE[6][78] ), 
        .D(\CACHE[7][78] ), .S0(n418), .S1(n450), .Y(n3257) );
  MXI4X1 U2504 ( .A(\CACHE[0][78] ), .B(\CACHE[1][78] ), .C(\CACHE[2][78] ), 
        .D(\CACHE[3][78] ), .S0(n418), .S1(n450), .Y(n3256) );
  MXI2X1 U2505 ( .A(n3258), .B(n3259), .S0(n469), .Y(N108) );
  MXI4X1 U2506 ( .A(\CACHE[4][79] ), .B(\CACHE[5][79] ), .C(\CACHE[6][79] ), 
        .D(\CACHE[7][79] ), .S0(n418), .S1(n450), .Y(n3259) );
  MXI4X1 U2507 ( .A(\CACHE[0][79] ), .B(\CACHE[1][79] ), .C(\CACHE[2][79] ), 
        .D(\CACHE[3][79] ), .S0(n418), .S1(n450), .Y(n3258) );
  MXI2X1 U2508 ( .A(n3260), .B(n3261), .S0(n470), .Y(N107) );
  MXI4X1 U2509 ( .A(\CACHE[4][80] ), .B(\CACHE[5][80] ), .C(\CACHE[6][80] ), 
        .D(\CACHE[7][80] ), .S0(n418), .S1(n450), .Y(n3261) );
  MXI4X1 U2510 ( .A(\CACHE[0][80] ), .B(\CACHE[1][80] ), .C(\CACHE[2][80] ), 
        .D(\CACHE[3][80] ), .S0(n418), .S1(n450), .Y(n3260) );
  MXI2X1 U2511 ( .A(n3262), .B(n3263), .S0(n468), .Y(N106) );
  MXI4X1 U2512 ( .A(\CACHE[4][81] ), .B(\CACHE[5][81] ), .C(\CACHE[6][81] ), 
        .D(\CACHE[7][81] ), .S0(n418), .S1(n450), .Y(n3263) );
  MXI4X1 U2513 ( .A(\CACHE[0][81] ), .B(\CACHE[1][81] ), .C(\CACHE[2][81] ), 
        .D(\CACHE[3][81] ), .S0(n418), .S1(n450), .Y(n3262) );
  MXI2X1 U2514 ( .A(n3264), .B(n3265), .S0(n467), .Y(N105) );
  MXI4X1 U2515 ( .A(\CACHE[4][82] ), .B(\CACHE[5][82] ), .C(\CACHE[6][82] ), 
        .D(\CACHE[7][82] ), .S0(n418), .S1(n450), .Y(n3265) );
  MXI4X1 U2516 ( .A(\CACHE[0][82] ), .B(\CACHE[1][82] ), .C(\CACHE[2][82] ), 
        .D(\CACHE[3][82] ), .S0(n418), .S1(n450), .Y(n3264) );
  MXI2X1 U2517 ( .A(n3266), .B(n3267), .S0(n468), .Y(N104) );
  MXI4X1 U2518 ( .A(\CACHE[4][83] ), .B(\CACHE[5][83] ), .C(\CACHE[6][83] ), 
        .D(\CACHE[7][83] ), .S0(n418), .S1(n450), .Y(n3267) );
  MXI4X1 U2519 ( .A(\CACHE[0][83] ), .B(\CACHE[1][83] ), .C(\CACHE[2][83] ), 
        .D(\CACHE[3][83] ), .S0(n418), .S1(n450), .Y(n3266) );
  MXI2X1 U2520 ( .A(n3268), .B(n3269), .S0(n473), .Y(N103) );
  MXI4X1 U2521 ( .A(\CACHE[4][84] ), .B(\CACHE[5][84] ), .C(\CACHE[6][84] ), 
        .D(\CACHE[7][84] ), .S0(n419), .S1(n451), .Y(n3269) );
  MXI4X1 U2522 ( .A(\CACHE[0][84] ), .B(\CACHE[1][84] ), .C(\CACHE[2][84] ), 
        .D(\CACHE[3][84] ), .S0(n419), .S1(n451), .Y(n3268) );
  MXI2X1 U2523 ( .A(n3270), .B(n3271), .S0(n473), .Y(N102) );
  MXI4X1 U2524 ( .A(\CACHE[4][85] ), .B(\CACHE[5][85] ), .C(\CACHE[6][85] ), 
        .D(\CACHE[7][85] ), .S0(n419), .S1(n451), .Y(n3271) );
  MXI4X1 U2525 ( .A(\CACHE[0][85] ), .B(\CACHE[1][85] ), .C(\CACHE[2][85] ), 
        .D(\CACHE[3][85] ), .S0(n419), .S1(n451), .Y(n3270) );
  MXI2X1 U2526 ( .A(n3272), .B(n3273), .S0(n473), .Y(N101) );
  MXI4X1 U2527 ( .A(\CACHE[4][86] ), .B(\CACHE[5][86] ), .C(\CACHE[6][86] ), 
        .D(\CACHE[7][86] ), .S0(n419), .S1(n451), .Y(n3273) );
  MXI4X1 U2528 ( .A(\CACHE[0][86] ), .B(\CACHE[1][86] ), .C(\CACHE[2][86] ), 
        .D(\CACHE[3][86] ), .S0(n419), .S1(n451), .Y(n3272) );
  MXI2X1 U2529 ( .A(n3274), .B(n3275), .S0(n473), .Y(N100) );
  MXI4X1 U2530 ( .A(\CACHE[4][87] ), .B(\CACHE[5][87] ), .C(\CACHE[6][87] ), 
        .D(\CACHE[7][87] ), .S0(n419), .S1(n451), .Y(n3275) );
  MXI4X1 U2531 ( .A(\CACHE[0][87] ), .B(\CACHE[1][87] ), .C(\CACHE[2][87] ), 
        .D(\CACHE[3][87] ), .S0(n419), .S1(n451), .Y(n3274) );
  MXI2X1 U2532 ( .A(n3276), .B(n3277), .S0(n471), .Y(N99) );
  MXI4X1 U2533 ( .A(\CACHE[4][88] ), .B(\CACHE[5][88] ), .C(\CACHE[6][88] ), 
        .D(\CACHE[7][88] ), .S0(n419), .S1(n451), .Y(n3277) );
  MXI4X1 U2534 ( .A(\CACHE[0][88] ), .B(\CACHE[1][88] ), .C(\CACHE[2][88] ), 
        .D(\CACHE[3][88] ), .S0(n419), .S1(n451), .Y(n3276) );
  MXI2X1 U2535 ( .A(n3278), .B(n3279), .S0(n464), .Y(N98) );
  MXI4X1 U2536 ( .A(\CACHE[4][89] ), .B(\CACHE[5][89] ), .C(\CACHE[6][89] ), 
        .D(\CACHE[7][89] ), .S0(n419), .S1(n451), .Y(n3279) );
  MXI4X1 U2537 ( .A(\CACHE[0][89] ), .B(\CACHE[1][89] ), .C(\CACHE[2][89] ), 
        .D(\CACHE[3][89] ), .S0(n419), .S1(n451), .Y(n3278) );
  MXI2X1 U2538 ( .A(n3280), .B(n3281), .S0(n465), .Y(N97) );
  MXI4X1 U2539 ( .A(\CACHE[4][90] ), .B(\CACHE[5][90] ), .C(\CACHE[6][90] ), 
        .D(\CACHE[7][90] ), .S0(n419), .S1(n452), .Y(n3281) );
  MXI4X1 U2540 ( .A(\CACHE[0][90] ), .B(\CACHE[1][90] ), .C(\CACHE[2][90] ), 
        .D(\CACHE[3][90] ), .S0(n419), .S1(n452), .Y(n3280) );
  MXI2X1 U2541 ( .A(n3282), .B(n3283), .S0(n466), .Y(N96) );
  MXI4X1 U2542 ( .A(\CACHE[4][91] ), .B(\CACHE[5][91] ), .C(\CACHE[6][91] ), 
        .D(\CACHE[7][91] ), .S0(n432), .S1(n452), .Y(n3283) );
  MXI4X1 U2543 ( .A(\CACHE[0][91] ), .B(\CACHE[1][91] ), .C(\CACHE[2][91] ), 
        .D(\CACHE[3][91] ), .S0(n436), .S1(n452), .Y(n3282) );
  MXI2X1 U2544 ( .A(n3284), .B(n3285), .S0(n469), .Y(N95) );
  MXI4X1 U2545 ( .A(\CACHE[4][92] ), .B(\CACHE[5][92] ), .C(\CACHE[6][92] ), 
        .D(\CACHE[7][92] ), .S0(n426), .S1(n452), .Y(n3285) );
  MXI4X1 U2546 ( .A(\CACHE[0][92] ), .B(\CACHE[1][92] ), .C(\CACHE[2][92] ), 
        .D(\CACHE[3][92] ), .S0(n433), .S1(n452), .Y(n3284) );
  MXI2X1 U2547 ( .A(n3286), .B(n3287), .S0(n470), .Y(N94) );
  MXI4X1 U2548 ( .A(\CACHE[4][93] ), .B(\CACHE[5][93] ), .C(\CACHE[6][93] ), 
        .D(\CACHE[7][93] ), .S0(n424), .S1(n452), .Y(n3287) );
  MXI4X1 U2549 ( .A(\CACHE[0][93] ), .B(\CACHE[1][93] ), .C(\CACHE[2][93] ), 
        .D(\CACHE[3][93] ), .S0(n429), .S1(n452), .Y(n3286) );
  MXI2X1 U2550 ( .A(n3288), .B(n3289), .S0(n465), .Y(N93) );
  MXI4X1 U2551 ( .A(\CACHE[4][94] ), .B(\CACHE[5][94] ), .C(\CACHE[6][94] ), 
        .D(\CACHE[7][94] ), .S0(n435), .S1(n452), .Y(n3289) );
  MXI4X1 U2552 ( .A(\CACHE[0][94] ), .B(\CACHE[1][94] ), .C(\CACHE[2][94] ), 
        .D(\CACHE[3][94] ), .S0(n425), .S1(n452), .Y(n3288) );
  MXI2X1 U2553 ( .A(n3290), .B(n3291), .S0(n467), .Y(N92) );
  MXI4X1 U2554 ( .A(\CACHE[4][95] ), .B(\CACHE[5][95] ), .C(\CACHE[6][95] ), 
        .D(\CACHE[7][95] ), .S0(n427), .S1(n452), .Y(n3291) );
  MXI4X1 U2555 ( .A(\CACHE[0][95] ), .B(\CACHE[1][95] ), .C(\CACHE[2][95] ), 
        .D(\CACHE[3][95] ), .S0(n428), .S1(n452), .Y(n3290) );
  NAND3BX1 U2556 ( .AN(n3408), .B(n3409), .C(n3410), .Y(proc_stall) );
  OAI221XL U2557 ( .A0(n3411), .A1(n3412), .B0(n3413), .B1(n3414), .C0(n3415), 
        .Y(proc_rdata[9]) );
  OAI221XL U2558 ( .A0(n3411), .A1(n3419), .B0(n3413), .B1(n3420), .C0(n3421), 
        .Y(proc_rdata[8]) );
  OAI221XL U2559 ( .A0(n3411), .A1(n3424), .B0(n3413), .B1(n3425), .C0(n3426), 
        .Y(proc_rdata[7]) );
  OAI221XL U2560 ( .A0(n3411), .A1(n3429), .B0(n3413), .B1(n3430), .C0(n3431), 
        .Y(proc_rdata[6]) );
  OAI221XL U2561 ( .A0(n3411), .A1(n3434), .B0(n3413), .B1(n3435), .C0(n3436), 
        .Y(proc_rdata[5]) );
  OAI221XL U2562 ( .A0(n3411), .A1(n3439), .B0(n3413), .B1(n3440), .C0(n3441), 
        .Y(proc_rdata[4]) );
  OAI221XL U2563 ( .A0(n3411), .A1(n3444), .B0(n3413), .B1(n3445), .C0(n3446), 
        .Y(proc_rdata[3]) );
  OAI221XL U2564 ( .A0(n3411), .A1(n3449), .B0(n3413), .B1(n3450), .C0(n3451), 
        .Y(proc_rdata[31]) );
  OAI221XL U2565 ( .A0(n3411), .A1(n3454), .B0(n3413), .B1(n3455), .C0(n3456), 
        .Y(proc_rdata[30]) );
  OAI221XL U2566 ( .A0(n3411), .A1(n3459), .B0(n3413), .B1(n3460), .C0(n3461), 
        .Y(proc_rdata[2]) );
  OAI221XL U2567 ( .A0(n3411), .A1(n3464), .B0(n3413), .B1(n3465), .C0(n3466), 
        .Y(proc_rdata[29]) );
  OAI221XL U2568 ( .A0(n3411), .A1(n3469), .B0(n3413), .B1(n3470), .C0(n3471), 
        .Y(proc_rdata[28]) );
  OAI221XL U2569 ( .A0(n3411), .A1(n3474), .B0(n3413), .B1(n3475), .C0(n3476), 
        .Y(proc_rdata[27]) );
  OAI221XL U2570 ( .A0(n3411), .A1(n3479), .B0(n3413), .B1(n3480), .C0(n3481), 
        .Y(proc_rdata[26]) );
  OAI221XL U2571 ( .A0(n3411), .A1(n3484), .B0(n3413), .B1(n3485), .C0(n3486), 
        .Y(proc_rdata[25]) );
  OAI221XL U2572 ( .A0(n3411), .A1(n3489), .B0(n3413), .B1(n3490), .C0(n3491), 
        .Y(proc_rdata[24]) );
  OAI221XL U2573 ( .A0(n3411), .A1(n3494), .B0(n3413), .B1(n3495), .C0(n3496), 
        .Y(proc_rdata[23]) );
  OAI221XL U2574 ( .A0(n3411), .A1(n3499), .B0(n3413), .B1(n3500), .C0(n3501), 
        .Y(proc_rdata[22]) );
  OAI221XL U2575 ( .A0(n3411), .A1(n3504), .B0(n3413), .B1(n3505), .C0(n3506), 
        .Y(proc_rdata[21]) );
  OAI221XL U2576 ( .A0(n3411), .A1(n3509), .B0(n3413), .B1(n3510), .C0(n3511), 
        .Y(proc_rdata[20]) );
  OAI221XL U2577 ( .A0(n3411), .A1(n3514), .B0(n3413), .B1(n3515), .C0(n3516), 
        .Y(proc_rdata[1]) );
  OAI221XL U2578 ( .A0(n3411), .A1(n3519), .B0(n3413), .B1(n3520), .C0(n3521), 
        .Y(proc_rdata[19]) );
  OAI221XL U2579 ( .A0(n3411), .A1(n3524), .B0(n3413), .B1(n3525), .C0(n3526), 
        .Y(proc_rdata[18]) );
  OAI221XL U2580 ( .A0(n3411), .A1(n3529), .B0(n3413), .B1(n3530), .C0(n3531), 
        .Y(proc_rdata[17]) );
  OAI221XL U2581 ( .A0(n3411), .A1(n3534), .B0(n3413), .B1(n3535), .C0(n3536), 
        .Y(proc_rdata[16]) );
  OAI221XL U2582 ( .A0(n3411), .A1(n3539), .B0(n3413), .B1(n3540), .C0(n3541), 
        .Y(proc_rdata[15]) );
  OAI221XL U2583 ( .A0(n3411), .A1(n3544), .B0(n3413), .B1(n3545), .C0(n3546), 
        .Y(proc_rdata[14]) );
  OAI221XL U2584 ( .A0(n3411), .A1(n3549), .B0(n3413), .B1(n3550), .C0(n3551), 
        .Y(proc_rdata[13]) );
  OAI221XL U2585 ( .A0(n3411), .A1(n3554), .B0(n3413), .B1(n3555), .C0(n3556), 
        .Y(proc_rdata[12]) );
  OAI221XL U2586 ( .A0(n3411), .A1(n3559), .B0(n3413), .B1(n3560), .C0(n3561), 
        .Y(proc_rdata[11]) );
  OAI221XL U2587 ( .A0(n3411), .A1(n3564), .B0(n3413), .B1(n3565), .C0(n3566), 
        .Y(proc_rdata[10]) );
  OAI221XL U2588 ( .A0(n3411), .A1(n3569), .B0(n3413), .B1(n3570), .C0(n3571), 
        .Y(proc_rdata[0]) );
  NOR3X1 U2589 ( .A(n462), .B(n437), .C(n475), .Y(n3578) );
  NOR3X1 U2590 ( .A(n462), .B(n436), .C(n474), .Y(n3733) );
  NOR3X1 U2591 ( .A(n438), .B(n460), .C(n474), .Y(n3734) );
  NOR3X1 U2592 ( .A(n423), .B(n460), .C(n475), .Y(n3735) );
  NOR3X1 U2593 ( .A(n437), .B(n472), .C(n461), .Y(n3736) );
  NOR3X1 U2594 ( .A(n421), .B(n472), .C(n461), .Y(n3737) );
  NOR3X1 U2595 ( .A(n460), .B(n473), .C(n439), .Y(n3738) );
  OAI31XL U2596 ( .A0(n3743), .A1(n3408), .A2(n3574), .B0(N34), .Y(n3741) );
  NAND3X1 U2597 ( .A(n3746), .B(n3742), .C(n3747), .Y(n3745) );
  OAI31XL U2598 ( .A0(n3751), .A1(n3575), .A2(n3576), .B0(n3752), .Y(n3750) );
  OAI31XL U2599 ( .A0(n3751), .A1(proc_addr[0]), .A2(n3576), .B0(n3752), .Y(
        n3755) );
  OAI31XL U2600 ( .A0(n3751), .A1(proc_addr[1]), .A2(n3575), .B0(n3752), .Y(
        n3758) );
  NOR3X1 U2601 ( .A(n444), .B(n473), .C(n436), .Y(n3739) );
  OAI31XL U2602 ( .A0(n3751), .A1(proc_addr[1]), .A2(proc_addr[0]), .B0(n3752), 
        .Y(n3761) );
  NAND2BX1 U2603 ( .AN(n3751), .B(n3742), .Y(n3752) );
  NOR2X1 U2604 ( .A(n3762), .B(n3763), .Y(n3740) );
  CLKINVX1 U2605 ( .A(n3766), .Y(n3765) );
  AOI21X1 U2606 ( .A0(n3764), .A1(N34), .B0(n3743), .Y(n3746) );
  OAI31XL U2607 ( .A0(n3410), .A1(N34), .A2(n3408), .B0(n3409), .Y(n3767) );
  CLKINVX1 U2608 ( .A(N178), .Y(n3416) );
  CLKINVX1 U2609 ( .A(N88), .Y(n3448) );
  CLKINVX1 U2610 ( .A(N89), .Y(n3463) );
  CLKINVX1 U2611 ( .A(N90), .Y(n3518) );
  CLKINVX1 U2612 ( .A(N91), .Y(n3573) );
  CLKINVX1 U2613 ( .A(N92), .Y(n3449) );
  CLKINVX1 U2614 ( .A(N93), .Y(n3454) );
  CLKINVX1 U2615 ( .A(N94), .Y(n3464) );
  CLKINVX1 U2616 ( .A(N95), .Y(n3469) );
  CLKINVX1 U2617 ( .A(N96), .Y(n3474) );
  CLKINVX1 U2618 ( .A(N97), .Y(n3479) );
  CLKINVX1 U2619 ( .A(N179), .Y(n3422) );
  CLKINVX1 U2620 ( .A(N98), .Y(n3484) );
  CLKINVX1 U2621 ( .A(N99), .Y(n3489) );
  CLKINVX1 U2622 ( .A(N100), .Y(n3494) );
  CLKINVX1 U2623 ( .A(N101), .Y(n3499) );
  CLKINVX1 U2624 ( .A(N102), .Y(n3504) );
  CLKINVX1 U2625 ( .A(N103), .Y(n3509) );
  CLKINVX1 U2626 ( .A(N104), .Y(n3519) );
  CLKINVX1 U2627 ( .A(N105), .Y(n3524) );
  CLKINVX1 U2628 ( .A(N106), .Y(n3529) );
  CLKINVX1 U2629 ( .A(N107), .Y(n3534) );
  CLKINVX1 U2630 ( .A(N180), .Y(n3427) );
  CLKINVX1 U2631 ( .A(N108), .Y(n3539) );
  CLKINVX1 U2632 ( .A(N109), .Y(n3544) );
  CLKINVX1 U2633 ( .A(N110), .Y(n3549) );
  CLKINVX1 U2634 ( .A(N111), .Y(n3554) );
  CLKINVX1 U2635 ( .A(N112), .Y(n3559) );
  CLKINVX1 U2636 ( .A(N113), .Y(n3564) );
  CLKINVX1 U2637 ( .A(N114), .Y(n3412) );
  CLKINVX1 U2638 ( .A(N115), .Y(n3419) );
  CLKINVX1 U2639 ( .A(N116), .Y(n3424) );
  CLKINVX1 U2640 ( .A(N117), .Y(n3429) );
  CLKINVX1 U2641 ( .A(N181), .Y(n3432) );
  CLKINVX1 U2642 ( .A(N118), .Y(n3434) );
  CLKINVX1 U2643 ( .A(N119), .Y(n3439) );
  CLKINVX1 U2644 ( .A(N120), .Y(n3444) );
  CLKINVX1 U2645 ( .A(N121), .Y(n3459) );
  CLKINVX1 U2646 ( .A(N122), .Y(n3514) );
  CLKINVX1 U2647 ( .A(N123), .Y(n3569) );
  CLKINVX1 U2648 ( .A(N124), .Y(n3450) );
  CLKINVX1 U2649 ( .A(N125), .Y(n3455) );
  CLKINVX1 U2650 ( .A(N126), .Y(n3465) );
  CLKINVX1 U2651 ( .A(N127), .Y(n3470) );
  CLKINVX1 U2652 ( .A(N182), .Y(n3437) );
  CLKINVX1 U2653 ( .A(N128), .Y(n3475) );
  CLKINVX1 U2654 ( .A(N129), .Y(n3480) );
  CLKINVX1 U2655 ( .A(N130), .Y(n3485) );
  CLKINVX1 U2656 ( .A(N131), .Y(n3490) );
  CLKINVX1 U2657 ( .A(N132), .Y(n3495) );
  CLKINVX1 U2658 ( .A(N133), .Y(n3500) );
  CLKINVX1 U2659 ( .A(N134), .Y(n3505) );
  CLKINVX1 U2660 ( .A(N135), .Y(n3510) );
  CLKINVX1 U2661 ( .A(N136), .Y(n3520) );
  CLKINVX1 U2662 ( .A(N137), .Y(n3525) );
  CLKINVX1 U2663 ( .A(N183), .Y(n3442) );
  CLKINVX1 U2664 ( .A(N138), .Y(n3530) );
  CLKINVX1 U2665 ( .A(N139), .Y(n3535) );
  CLKINVX1 U2666 ( .A(N140), .Y(n3540) );
  CLKINVX1 U2667 ( .A(N141), .Y(n3545) );
  CLKINVX1 U2668 ( .A(N142), .Y(n3550) );
  CLKINVX1 U2669 ( .A(N143), .Y(n3555) );
  CLKINVX1 U2670 ( .A(N144), .Y(n3560) );
  CLKINVX1 U2671 ( .A(N145), .Y(n3565) );
  CLKINVX1 U2672 ( .A(N146), .Y(n3414) );
  CLKINVX1 U2673 ( .A(N147), .Y(n3420) );
  CLKINVX1 U2674 ( .A(N184), .Y(n3447) );
  CLKINVX1 U2675 ( .A(N148), .Y(n3425) );
  CLKINVX1 U2676 ( .A(N149), .Y(n3430) );
  CLKINVX1 U2677 ( .A(N150), .Y(n3435) );
  CLKINVX1 U2678 ( .A(N151), .Y(n3440) );
  CLKINVX1 U2679 ( .A(N152), .Y(n3445) );
  CLKINVX1 U2680 ( .A(N153), .Y(n3460) );
  CLKINVX1 U2681 ( .A(N154), .Y(n3515) );
  CLKINVX1 U2682 ( .A(N155), .Y(n3570) );
  CLKINVX1 U2683 ( .A(N156), .Y(n3452) );
  CLKINVX1 U2684 ( .A(N157), .Y(n3457) );
  CLKINVX1 U2685 ( .A(N185), .Y(n3462) );
  CLKINVX1 U2686 ( .A(N158), .Y(n3467) );
  CLKINVX1 U2687 ( .A(N159), .Y(n3472) );
  CLKINVX1 U2688 ( .A(N160), .Y(n3477) );
  CLKINVX1 U2689 ( .A(N161), .Y(n3482) );
  CLKINVX1 U2690 ( .A(N162), .Y(n3487) );
  CLKINVX1 U2691 ( .A(N163), .Y(n3492) );
  CLKINVX1 U2692 ( .A(N164), .Y(n3497) );
  CLKINVX1 U2693 ( .A(N165), .Y(n3502) );
  CLKINVX1 U2694 ( .A(N166), .Y(n3507) );
  CLKINVX1 U2695 ( .A(N167), .Y(n3512) );
  CLKINVX1 U2696 ( .A(N186), .Y(n3517) );
  CLKINVX1 U2697 ( .A(N168), .Y(n3522) );
  CLKINVX1 U2698 ( .A(N169), .Y(n3527) );
  CLKINVX1 U2699 ( .A(N170), .Y(n3532) );
  CLKINVX1 U2700 ( .A(N171), .Y(n3537) );
  CLKINVX1 U2701 ( .A(N172), .Y(n3542) );
  CLKINVX1 U2702 ( .A(N173), .Y(n3547) );
  CLKINVX1 U2703 ( .A(N174), .Y(n3552) );
  CLKINVX1 U2704 ( .A(N175), .Y(n3557) );
  CLKINVX1 U2705 ( .A(N60), .Y(n3453) );
  CLKINVX1 U2706 ( .A(N61), .Y(n3458) );
  CLKINVX1 U2707 ( .A(N62), .Y(n3468) );
  CLKINVX1 U2708 ( .A(N63), .Y(n3473) );
  CLKINVX1 U2709 ( .A(N64), .Y(n3478) );
  CLKINVX1 U2710 ( .A(N65), .Y(n3483) );
  CLKINVX1 U2711 ( .A(N66), .Y(n3488) );
  CLKINVX1 U2712 ( .A(N67), .Y(n3493) );
  CLKINVX1 U2713 ( .A(N176), .Y(n3562) );
  CLKINVX1 U2714 ( .A(N68), .Y(n3498) );
  CLKINVX1 U2715 ( .A(N69), .Y(n3503) );
  CLKINVX1 U2716 ( .A(N70), .Y(n3508) );
  CLKINVX1 U2717 ( .A(N71), .Y(n3513) );
  CLKINVX1 U2718 ( .A(N72), .Y(n3523) );
  CLKINVX1 U2719 ( .A(N73), .Y(n3528) );
  CLKINVX1 U2720 ( .A(N74), .Y(n3533) );
  CLKINVX1 U2721 ( .A(N75), .Y(n3538) );
  CLKINVX1 U2722 ( .A(N76), .Y(n3543) );
  CLKINVX1 U2723 ( .A(N77), .Y(n3548) );
  CLKINVX1 U2724 ( .A(N177), .Y(n3567) );
  CLKINVX1 U2725 ( .A(N78), .Y(n3553) );
  CLKINVX1 U2726 ( .A(N79), .Y(n3558) );
  CLKINVX1 U2727 ( .A(N80), .Y(n3563) );
  CLKINVX1 U2728 ( .A(N81), .Y(n3568) );
  CLKINVX1 U2729 ( .A(N82), .Y(n3418) );
  CLKINVX1 U2730 ( .A(N83), .Y(n3423) );
  CLKINVX1 U2731 ( .A(N84), .Y(n3428) );
  CLKINVX1 U2732 ( .A(N85), .Y(n3433) );
  CLKINVX1 U2733 ( .A(N86), .Y(n3438) );
  CLKINVX1 U2734 ( .A(N87), .Y(n3443) );
  CLKINVX1 U2735 ( .A(N187), .Y(n3572) );
  NOR2X1 U2736 ( .A(n413), .B(mem_read), .Y(n3768) );
  NOR3BXL U2737 ( .AN(n3769), .B(n3408), .C(mem_ready), .Y(n3804) );
  NOR2X1 U2738 ( .A(proc_read), .B(proc_write), .Y(n3408) );
  OAI21XL U2739 ( .A0(N34), .A1(n3410), .B0(n3409), .Y(n3769) );
  NAND2BX1 U2740 ( .AN(N33), .B(proc_read), .Y(n3409) );
  CLKINVX1 U2741 ( .A(n3763), .Y(n3410) );
  CLKINVX1 U2742 ( .A(mem_ready), .Y(n3743) );
  NAND4X1 U2743 ( .A(n3771), .B(n3772), .C(n3773), .D(n3774), .Y(n3763) );
  NOR4X1 U2744 ( .A(n3775), .B(n3776), .C(n3777), .D(n3778), .Y(n3774) );
  NAND4X1 U2745 ( .A(n3779), .B(n3780), .C(n3781), .D(n3782), .Y(n3775) );
  NOR4X1 U2746 ( .A(n3783), .B(n3784), .C(n3785), .D(n3786), .Y(n3773) );
  NAND3X1 U2747 ( .A(n3787), .B(n3788), .C(n3789), .Y(n3783) );
  NOR4X1 U2748 ( .A(n3790), .B(n3791), .C(n3792), .D(n3793), .Y(n3772) );
  NAND3X1 U2749 ( .A(n3794), .B(n3795), .C(n3796), .Y(n3790) );
  NOR4X1 U2750 ( .A(n3797), .B(n3798), .C(n3799), .D(n3800), .Y(n3771) );
  NAND3X1 U2751 ( .A(n3801), .B(n3802), .C(n3803), .Y(n3797) );
  NAND2X1 U2752 ( .A(n3762), .B(n3766), .Y(n3770) );
  NAND2X1 U2753 ( .A(N33), .B(proc_read), .Y(n3766) );
  CLKINVX1 U2754 ( .A(proc_read), .Y(n3764) );
endmodule


module cache_1 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N30, N31, N32, n6281, \CACHE[7][154] , \CACHE[7][153] ,
         \CACHE[7][152] , \CACHE[7][151] , \CACHE[7][150] , \CACHE[7][149] ,
         \CACHE[7][148] , \CACHE[7][147] , \CACHE[7][146] , \CACHE[7][145] ,
         \CACHE[7][144] , \CACHE[7][143] , \CACHE[7][142] , \CACHE[7][141] ,
         \CACHE[7][140] , \CACHE[7][139] , \CACHE[7][138] , \CACHE[7][137] ,
         \CACHE[7][136] , \CACHE[7][135] , \CACHE[7][134] , \CACHE[7][133] ,
         \CACHE[7][132] , \CACHE[7][131] , \CACHE[7][130] , \CACHE[7][129] ,
         \CACHE[7][128] , \CACHE[7][127] , \CACHE[7][126] , \CACHE[7][125] ,
         \CACHE[7][124] , \CACHE[7][123] , \CACHE[7][122] , \CACHE[7][121] ,
         \CACHE[7][120] , \CACHE[7][119] , \CACHE[7][118] , \CACHE[7][117] ,
         \CACHE[7][116] , \CACHE[7][115] , \CACHE[7][114] , \CACHE[7][113] ,
         \CACHE[7][112] , \CACHE[7][111] , \CACHE[7][110] , \CACHE[7][109] ,
         \CACHE[7][108] , \CACHE[7][107] , \CACHE[7][106] , \CACHE[7][105] ,
         \CACHE[7][104] , \CACHE[7][103] , \CACHE[7][102] , \CACHE[7][101] ,
         \CACHE[7][100] , \CACHE[7][99] , \CACHE[7][98] , \CACHE[7][97] ,
         \CACHE[7][96] , \CACHE[7][95] , \CACHE[7][94] , \CACHE[7][93] ,
         \CACHE[7][92] , \CACHE[7][91] , \CACHE[7][90] , \CACHE[7][89] ,
         \CACHE[7][88] , \CACHE[7][87] , \CACHE[7][86] , \CACHE[7][85] ,
         \CACHE[7][84] , \CACHE[7][83] , \CACHE[7][82] , \CACHE[7][81] ,
         \CACHE[7][80] , \CACHE[7][79] , \CACHE[7][78] , \CACHE[7][77] ,
         \CACHE[7][76] , \CACHE[7][75] , \CACHE[7][74] , \CACHE[7][73] ,
         \CACHE[7][72] , \CACHE[7][71] , \CACHE[7][70] , \CACHE[7][69] ,
         \CACHE[7][68] , \CACHE[7][67] , \CACHE[7][66] , \CACHE[7][65] ,
         \CACHE[7][64] , \CACHE[7][63] , \CACHE[7][62] , \CACHE[7][61] ,
         \CACHE[7][60] , \CACHE[7][59] , \CACHE[7][58] , \CACHE[7][57] ,
         \CACHE[7][56] , \CACHE[7][55] , \CACHE[7][54] , \CACHE[7][53] ,
         \CACHE[7][52] , \CACHE[7][51] , \CACHE[7][50] , \CACHE[7][49] ,
         \CACHE[7][48] , \CACHE[7][47] , \CACHE[7][46] , \CACHE[7][45] ,
         \CACHE[7][44] , \CACHE[7][43] , \CACHE[7][42] , \CACHE[7][41] ,
         \CACHE[7][40] , \CACHE[7][39] , \CACHE[7][38] , \CACHE[7][37] ,
         \CACHE[7][36] , \CACHE[7][35] , \CACHE[7][34] , \CACHE[7][33] ,
         \CACHE[7][32] , \CACHE[7][31] , \CACHE[7][30] , \CACHE[7][29] ,
         \CACHE[7][28] , \CACHE[7][27] , \CACHE[7][26] , \CACHE[7][25] ,
         \CACHE[7][24] , \CACHE[7][23] , \CACHE[7][22] , \CACHE[7][21] ,
         \CACHE[7][20] , \CACHE[7][19] , \CACHE[7][18] , \CACHE[7][17] ,
         \CACHE[7][16] , \CACHE[7][15] , \CACHE[7][14] , \CACHE[7][13] ,
         \CACHE[7][12] , \CACHE[7][11] , \CACHE[7][10] , \CACHE[7][9] ,
         \CACHE[7][8] , \CACHE[7][7] , \CACHE[7][6] , \CACHE[7][5] ,
         \CACHE[7][4] , \CACHE[7][3] , \CACHE[7][2] , \CACHE[7][1] ,
         \CACHE[7][0] , \CACHE[6][154] , \CACHE[6][153] , \CACHE[6][152] ,
         \CACHE[6][151] , \CACHE[6][150] , \CACHE[6][149] , \CACHE[6][148] ,
         \CACHE[6][147] , \CACHE[6][146] , \CACHE[6][145] , \CACHE[6][144] ,
         \CACHE[6][143] , \CACHE[6][142] , \CACHE[6][141] , \CACHE[6][140] ,
         \CACHE[6][139] , \CACHE[6][138] , \CACHE[6][137] , \CACHE[6][136] ,
         \CACHE[6][135] , \CACHE[6][134] , \CACHE[6][133] , \CACHE[6][132] ,
         \CACHE[6][131] , \CACHE[6][130] , \CACHE[6][129] , \CACHE[6][128] ,
         \CACHE[6][127] , \CACHE[6][126] , \CACHE[6][125] , \CACHE[6][124] ,
         \CACHE[6][123] , \CACHE[6][122] , \CACHE[6][121] , \CACHE[6][120] ,
         \CACHE[6][119] , \CACHE[6][118] , \CACHE[6][117] , \CACHE[6][116] ,
         \CACHE[6][115] , \CACHE[6][114] , \CACHE[6][113] , \CACHE[6][112] ,
         \CACHE[6][111] , \CACHE[6][110] , \CACHE[6][109] , \CACHE[6][108] ,
         \CACHE[6][107] , \CACHE[6][106] , \CACHE[6][105] , \CACHE[6][104] ,
         \CACHE[6][103] , \CACHE[6][102] , \CACHE[6][101] , \CACHE[6][100] ,
         \CACHE[6][99] , \CACHE[6][98] , \CACHE[6][97] , \CACHE[6][96] ,
         \CACHE[6][95] , \CACHE[6][94] , \CACHE[6][93] , \CACHE[6][92] ,
         \CACHE[6][91] , \CACHE[6][90] , \CACHE[6][89] , \CACHE[6][88] ,
         \CACHE[6][87] , \CACHE[6][86] , \CACHE[6][85] , \CACHE[6][84] ,
         \CACHE[6][83] , \CACHE[6][82] , \CACHE[6][81] , \CACHE[6][80] ,
         \CACHE[6][79] , \CACHE[6][78] , \CACHE[6][77] , \CACHE[6][76] ,
         \CACHE[6][75] , \CACHE[6][74] , \CACHE[6][73] , \CACHE[6][72] ,
         \CACHE[6][71] , \CACHE[6][70] , \CACHE[6][69] , \CACHE[6][68] ,
         \CACHE[6][67] , \CACHE[6][66] , \CACHE[6][65] , \CACHE[6][64] ,
         \CACHE[6][63] , \CACHE[6][62] , \CACHE[6][61] , \CACHE[6][60] ,
         \CACHE[6][59] , \CACHE[6][58] , \CACHE[6][57] , \CACHE[6][56] ,
         \CACHE[6][55] , \CACHE[6][54] , \CACHE[6][53] , \CACHE[6][52] ,
         \CACHE[6][51] , \CACHE[6][50] , \CACHE[6][49] , \CACHE[6][48] ,
         \CACHE[6][47] , \CACHE[6][46] , \CACHE[6][45] , \CACHE[6][44] ,
         \CACHE[6][43] , \CACHE[6][42] , \CACHE[6][41] , \CACHE[6][40] ,
         \CACHE[6][39] , \CACHE[6][38] , \CACHE[6][37] , \CACHE[6][36] ,
         \CACHE[6][35] , \CACHE[6][34] , \CACHE[6][33] , \CACHE[6][32] ,
         \CACHE[6][31] , \CACHE[6][30] , \CACHE[6][29] , \CACHE[6][28] ,
         \CACHE[6][27] , \CACHE[6][26] , \CACHE[6][25] , \CACHE[6][24] ,
         \CACHE[6][23] , \CACHE[6][22] , \CACHE[6][21] , \CACHE[6][20] ,
         \CACHE[6][19] , \CACHE[6][18] , \CACHE[6][17] , \CACHE[6][16] ,
         \CACHE[6][15] , \CACHE[6][14] , \CACHE[6][13] , \CACHE[6][12] ,
         \CACHE[6][11] , \CACHE[6][10] , \CACHE[6][9] , \CACHE[6][8] ,
         \CACHE[6][7] , \CACHE[6][6] , \CACHE[6][5] , \CACHE[6][4] ,
         \CACHE[6][3] , \CACHE[6][2] , \CACHE[6][1] , \CACHE[6][0] ,
         \CACHE[5][154] , \CACHE[5][153] , \CACHE[5][152] , \CACHE[5][151] ,
         \CACHE[5][150] , \CACHE[5][149] , \CACHE[5][148] , \CACHE[5][147] ,
         \CACHE[5][146] , \CACHE[5][145] , \CACHE[5][144] , \CACHE[5][143] ,
         \CACHE[5][142] , \CACHE[5][141] , \CACHE[5][140] , \CACHE[5][139] ,
         \CACHE[5][138] , \CACHE[5][137] , \CACHE[5][136] , \CACHE[5][135] ,
         \CACHE[5][134] , \CACHE[5][133] , \CACHE[5][132] , \CACHE[5][131] ,
         \CACHE[5][130] , \CACHE[5][129] , \CACHE[5][128] , \CACHE[5][127] ,
         \CACHE[5][126] , \CACHE[5][125] , \CACHE[5][124] , \CACHE[5][123] ,
         \CACHE[5][122] , \CACHE[5][121] , \CACHE[5][120] , \CACHE[5][119] ,
         \CACHE[5][118] , \CACHE[5][117] , \CACHE[5][116] , \CACHE[5][115] ,
         \CACHE[5][114] , \CACHE[5][113] , \CACHE[5][112] , \CACHE[5][111] ,
         \CACHE[5][110] , \CACHE[5][109] , \CACHE[5][108] , \CACHE[5][107] ,
         \CACHE[5][106] , \CACHE[5][105] , \CACHE[5][104] , \CACHE[5][103] ,
         \CACHE[5][102] , \CACHE[5][101] , \CACHE[5][100] , \CACHE[5][99] ,
         \CACHE[5][98] , \CACHE[5][97] , \CACHE[5][96] , \CACHE[5][95] ,
         \CACHE[5][94] , \CACHE[5][93] , \CACHE[5][92] , \CACHE[5][91] ,
         \CACHE[5][90] , \CACHE[5][89] , \CACHE[5][88] , \CACHE[5][87] ,
         \CACHE[5][86] , \CACHE[5][85] , \CACHE[5][84] , \CACHE[5][83] ,
         \CACHE[5][82] , \CACHE[5][81] , \CACHE[5][80] , \CACHE[5][79] ,
         \CACHE[5][78] , \CACHE[5][77] , \CACHE[5][76] , \CACHE[5][75] ,
         \CACHE[5][74] , \CACHE[5][73] , \CACHE[5][72] , \CACHE[5][71] ,
         \CACHE[5][70] , \CACHE[5][69] , \CACHE[5][68] , \CACHE[5][67] ,
         \CACHE[5][66] , \CACHE[5][65] , \CACHE[5][64] , \CACHE[5][63] ,
         \CACHE[5][62] , \CACHE[5][61] , \CACHE[5][60] , \CACHE[5][59] ,
         \CACHE[5][58] , \CACHE[5][57] , \CACHE[5][56] , \CACHE[5][55] ,
         \CACHE[5][54] , \CACHE[5][53] , \CACHE[5][52] , \CACHE[5][51] ,
         \CACHE[5][50] , \CACHE[5][49] , \CACHE[5][48] , \CACHE[5][47] ,
         \CACHE[5][46] , \CACHE[5][45] , \CACHE[5][44] , \CACHE[5][43] ,
         \CACHE[5][42] , \CACHE[5][41] , \CACHE[5][40] , \CACHE[5][39] ,
         \CACHE[5][38] , \CACHE[5][37] , \CACHE[5][36] , \CACHE[5][35] ,
         \CACHE[5][34] , \CACHE[5][33] , \CACHE[5][32] , \CACHE[5][31] ,
         \CACHE[5][30] , \CACHE[5][29] , \CACHE[5][28] , \CACHE[5][27] ,
         \CACHE[5][26] , \CACHE[5][25] , \CACHE[5][24] , \CACHE[5][23] ,
         \CACHE[5][22] , \CACHE[5][21] , \CACHE[5][20] , \CACHE[5][19] ,
         \CACHE[5][18] , \CACHE[5][17] , \CACHE[5][16] , \CACHE[5][15] ,
         \CACHE[5][14] , \CACHE[5][13] , \CACHE[5][12] , \CACHE[5][11] ,
         \CACHE[5][10] , \CACHE[5][9] , \CACHE[5][8] , \CACHE[5][7] ,
         \CACHE[5][6] , \CACHE[5][5] , \CACHE[5][4] , \CACHE[5][3] ,
         \CACHE[5][2] , \CACHE[5][1] , \CACHE[5][0] , \CACHE[4][154] ,
         \CACHE[4][153] , \CACHE[4][152] , \CACHE[4][151] , \CACHE[4][150] ,
         \CACHE[4][149] , \CACHE[4][148] , \CACHE[4][147] , \CACHE[4][146] ,
         \CACHE[4][145] , \CACHE[4][144] , \CACHE[4][143] , \CACHE[4][142] ,
         \CACHE[4][141] , \CACHE[4][140] , \CACHE[4][139] , \CACHE[4][138] ,
         \CACHE[4][137] , \CACHE[4][136] , \CACHE[4][135] , \CACHE[4][134] ,
         \CACHE[4][133] , \CACHE[4][132] , \CACHE[4][131] , \CACHE[4][130] ,
         \CACHE[4][129] , \CACHE[4][128] , \CACHE[4][127] , \CACHE[4][126] ,
         \CACHE[4][125] , \CACHE[4][124] , \CACHE[4][123] , \CACHE[4][122] ,
         \CACHE[4][121] , \CACHE[4][120] , \CACHE[4][119] , \CACHE[4][118] ,
         \CACHE[4][117] , \CACHE[4][116] , \CACHE[4][115] , \CACHE[4][114] ,
         \CACHE[4][113] , \CACHE[4][112] , \CACHE[4][111] , \CACHE[4][110] ,
         \CACHE[4][109] , \CACHE[4][108] , \CACHE[4][107] , \CACHE[4][106] ,
         \CACHE[4][105] , \CACHE[4][104] , \CACHE[4][103] , \CACHE[4][102] ,
         \CACHE[4][101] , \CACHE[4][100] , \CACHE[4][99] , \CACHE[4][98] ,
         \CACHE[4][97] , \CACHE[4][96] , \CACHE[4][95] , \CACHE[4][94] ,
         \CACHE[4][93] , \CACHE[4][92] , \CACHE[4][91] , \CACHE[4][90] ,
         \CACHE[4][89] , \CACHE[4][88] , \CACHE[4][87] , \CACHE[4][86] ,
         \CACHE[4][85] , \CACHE[4][84] , \CACHE[4][83] , \CACHE[4][82] ,
         \CACHE[4][81] , \CACHE[4][80] , \CACHE[4][79] , \CACHE[4][78] ,
         \CACHE[4][77] , \CACHE[4][76] , \CACHE[4][75] , \CACHE[4][74] ,
         \CACHE[4][73] , \CACHE[4][72] , \CACHE[4][71] , \CACHE[4][70] ,
         \CACHE[4][69] , \CACHE[4][68] , \CACHE[4][67] , \CACHE[4][66] ,
         \CACHE[4][65] , \CACHE[4][64] , \CACHE[4][63] , \CACHE[4][62] ,
         \CACHE[4][61] , \CACHE[4][60] , \CACHE[4][59] , \CACHE[4][58] ,
         \CACHE[4][57] , \CACHE[4][56] , \CACHE[4][55] , \CACHE[4][54] ,
         \CACHE[4][53] , \CACHE[4][52] , \CACHE[4][51] , \CACHE[4][50] ,
         \CACHE[4][49] , \CACHE[4][48] , \CACHE[4][47] , \CACHE[4][46] ,
         \CACHE[4][45] , \CACHE[4][44] , \CACHE[4][43] , \CACHE[4][42] ,
         \CACHE[4][41] , \CACHE[4][40] , \CACHE[4][39] , \CACHE[4][38] ,
         \CACHE[4][37] , \CACHE[4][36] , \CACHE[4][35] , \CACHE[4][34] ,
         \CACHE[4][33] , \CACHE[4][32] , \CACHE[4][31] , \CACHE[4][30] ,
         \CACHE[4][29] , \CACHE[4][28] , \CACHE[4][27] , \CACHE[4][26] ,
         \CACHE[4][25] , \CACHE[4][24] , \CACHE[4][23] , \CACHE[4][22] ,
         \CACHE[4][21] , \CACHE[4][20] , \CACHE[4][19] , \CACHE[4][18] ,
         \CACHE[4][17] , \CACHE[4][16] , \CACHE[4][15] , \CACHE[4][14] ,
         \CACHE[4][13] , \CACHE[4][12] , \CACHE[4][11] , \CACHE[4][10] ,
         \CACHE[4][9] , \CACHE[4][8] , \CACHE[4][7] , \CACHE[4][6] ,
         \CACHE[4][5] , \CACHE[4][4] , \CACHE[4][3] , \CACHE[4][2] ,
         \CACHE[4][1] , \CACHE[4][0] , \CACHE[3][154] , \CACHE[3][153] ,
         \CACHE[3][152] , \CACHE[3][151] , \CACHE[3][150] , \CACHE[3][149] ,
         \CACHE[3][148] , \CACHE[3][147] , \CACHE[3][146] , \CACHE[3][145] ,
         \CACHE[3][144] , \CACHE[3][143] , \CACHE[3][142] , \CACHE[3][141] ,
         \CACHE[3][140] , \CACHE[3][139] , \CACHE[3][138] , \CACHE[3][137] ,
         \CACHE[3][136] , \CACHE[3][135] , \CACHE[3][134] , \CACHE[3][133] ,
         \CACHE[3][132] , \CACHE[3][131] , \CACHE[3][130] , \CACHE[3][129] ,
         \CACHE[3][128] , \CACHE[3][127] , \CACHE[3][126] , \CACHE[3][125] ,
         \CACHE[3][124] , \CACHE[3][123] , \CACHE[3][122] , \CACHE[3][121] ,
         \CACHE[3][120] , \CACHE[3][119] , \CACHE[3][118] , \CACHE[3][117] ,
         \CACHE[3][116] , \CACHE[3][115] , \CACHE[3][114] , \CACHE[3][113] ,
         \CACHE[3][112] , \CACHE[3][111] , \CACHE[3][110] , \CACHE[3][109] ,
         \CACHE[3][108] , \CACHE[3][107] , \CACHE[3][106] , \CACHE[3][105] ,
         \CACHE[3][104] , \CACHE[3][103] , \CACHE[3][102] , \CACHE[3][101] ,
         \CACHE[3][100] , \CACHE[3][99] , \CACHE[3][98] , \CACHE[3][97] ,
         \CACHE[3][96] , \CACHE[3][95] , \CACHE[3][94] , \CACHE[3][93] ,
         \CACHE[3][92] , \CACHE[3][91] , \CACHE[3][90] , \CACHE[3][89] ,
         \CACHE[3][88] , \CACHE[3][87] , \CACHE[3][86] , \CACHE[3][85] ,
         \CACHE[3][84] , \CACHE[3][83] , \CACHE[3][82] , \CACHE[3][81] ,
         \CACHE[3][80] , \CACHE[3][79] , \CACHE[3][78] , \CACHE[3][77] ,
         \CACHE[3][76] , \CACHE[3][75] , \CACHE[3][74] , \CACHE[3][73] ,
         \CACHE[3][72] , \CACHE[3][71] , \CACHE[3][70] , \CACHE[3][69] ,
         \CACHE[3][68] , \CACHE[3][67] , \CACHE[3][66] , \CACHE[3][65] ,
         \CACHE[3][64] , \CACHE[3][63] , \CACHE[3][62] , \CACHE[3][61] ,
         \CACHE[3][60] , \CACHE[3][59] , \CACHE[3][58] , \CACHE[3][57] ,
         \CACHE[3][56] , \CACHE[3][55] , \CACHE[3][54] , \CACHE[3][53] ,
         \CACHE[3][52] , \CACHE[3][51] , \CACHE[3][50] , \CACHE[3][49] ,
         \CACHE[3][48] , \CACHE[3][47] , \CACHE[3][46] , \CACHE[3][45] ,
         \CACHE[3][44] , \CACHE[3][43] , \CACHE[3][42] , \CACHE[3][41] ,
         \CACHE[3][40] , \CACHE[3][39] , \CACHE[3][38] , \CACHE[3][37] ,
         \CACHE[3][36] , \CACHE[3][35] , \CACHE[3][34] , \CACHE[3][33] ,
         \CACHE[3][32] , \CACHE[3][31] , \CACHE[3][30] , \CACHE[3][29] ,
         \CACHE[3][28] , \CACHE[3][27] , \CACHE[3][26] , \CACHE[3][25] ,
         \CACHE[3][24] , \CACHE[3][23] , \CACHE[3][22] , \CACHE[3][21] ,
         \CACHE[3][20] , \CACHE[3][19] , \CACHE[3][18] , \CACHE[3][17] ,
         \CACHE[3][16] , \CACHE[3][15] , \CACHE[3][14] , \CACHE[3][13] ,
         \CACHE[3][12] , \CACHE[3][11] , \CACHE[3][10] , \CACHE[3][9] ,
         \CACHE[3][8] , \CACHE[3][7] , \CACHE[3][6] , \CACHE[3][5] ,
         \CACHE[3][4] , \CACHE[3][3] , \CACHE[3][2] , \CACHE[3][1] ,
         \CACHE[3][0] , \CACHE[2][154] , \CACHE[2][153] , \CACHE[2][152] ,
         \CACHE[2][151] , \CACHE[2][150] , \CACHE[2][149] , \CACHE[2][148] ,
         \CACHE[2][147] , \CACHE[2][146] , \CACHE[2][145] , \CACHE[2][144] ,
         \CACHE[2][143] , \CACHE[2][142] , \CACHE[2][141] , \CACHE[2][140] ,
         \CACHE[2][139] , \CACHE[2][138] , \CACHE[2][137] , \CACHE[2][136] ,
         \CACHE[2][135] , \CACHE[2][134] , \CACHE[2][133] , \CACHE[2][132] ,
         \CACHE[2][131] , \CACHE[2][130] , \CACHE[2][129] , \CACHE[2][128] ,
         \CACHE[2][127] , \CACHE[2][126] , \CACHE[2][125] , \CACHE[2][124] ,
         \CACHE[2][123] , \CACHE[2][122] , \CACHE[2][121] , \CACHE[2][120] ,
         \CACHE[2][119] , \CACHE[2][118] , \CACHE[2][117] , \CACHE[2][116] ,
         \CACHE[2][115] , \CACHE[2][114] , \CACHE[2][113] , \CACHE[2][112] ,
         \CACHE[2][111] , \CACHE[2][110] , \CACHE[2][109] , \CACHE[2][108] ,
         \CACHE[2][107] , \CACHE[2][106] , \CACHE[2][105] , \CACHE[2][104] ,
         \CACHE[2][103] , \CACHE[2][102] , \CACHE[2][101] , \CACHE[2][100] ,
         \CACHE[2][99] , \CACHE[2][98] , \CACHE[2][97] , \CACHE[2][96] ,
         \CACHE[2][95] , \CACHE[2][94] , \CACHE[2][93] , \CACHE[2][92] ,
         \CACHE[2][91] , \CACHE[2][90] , \CACHE[2][89] , \CACHE[2][88] ,
         \CACHE[2][87] , \CACHE[2][86] , \CACHE[2][85] , \CACHE[2][84] ,
         \CACHE[2][83] , \CACHE[2][82] , \CACHE[2][81] , \CACHE[2][80] ,
         \CACHE[2][79] , \CACHE[2][78] , \CACHE[2][77] , \CACHE[2][76] ,
         \CACHE[2][75] , \CACHE[2][74] , \CACHE[2][73] , \CACHE[2][72] ,
         \CACHE[2][71] , \CACHE[2][70] , \CACHE[2][69] , \CACHE[2][68] ,
         \CACHE[2][67] , \CACHE[2][66] , \CACHE[2][65] , \CACHE[2][64] ,
         \CACHE[2][63] , \CACHE[2][62] , \CACHE[2][61] , \CACHE[2][60] ,
         \CACHE[2][59] , \CACHE[2][58] , \CACHE[2][57] , \CACHE[2][56] ,
         \CACHE[2][55] , \CACHE[2][54] , \CACHE[2][53] , \CACHE[2][52] ,
         \CACHE[2][51] , \CACHE[2][50] , \CACHE[2][49] , \CACHE[2][48] ,
         \CACHE[2][47] , \CACHE[2][46] , \CACHE[2][45] , \CACHE[2][44] ,
         \CACHE[2][43] , \CACHE[2][42] , \CACHE[2][41] , \CACHE[2][40] ,
         \CACHE[2][39] , \CACHE[2][38] , \CACHE[2][37] , \CACHE[2][36] ,
         \CACHE[2][35] , \CACHE[2][34] , \CACHE[2][33] , \CACHE[2][32] ,
         \CACHE[2][31] , \CACHE[2][30] , \CACHE[2][29] , \CACHE[2][28] ,
         \CACHE[2][27] , \CACHE[2][26] , \CACHE[2][25] , \CACHE[2][24] ,
         \CACHE[2][23] , \CACHE[2][22] , \CACHE[2][21] , \CACHE[2][20] ,
         \CACHE[2][19] , \CACHE[2][18] , \CACHE[2][17] , \CACHE[2][16] ,
         \CACHE[2][15] , \CACHE[2][14] , \CACHE[2][13] , \CACHE[2][12] ,
         \CACHE[2][11] , \CACHE[2][10] , \CACHE[2][9] , \CACHE[2][8] ,
         \CACHE[2][7] , \CACHE[2][6] , \CACHE[2][5] , \CACHE[2][4] ,
         \CACHE[2][3] , \CACHE[2][2] , \CACHE[2][1] , \CACHE[2][0] ,
         \CACHE[1][154] , \CACHE[1][153] , \CACHE[1][152] , \CACHE[1][151] ,
         \CACHE[1][150] , \CACHE[1][149] , \CACHE[1][148] , \CACHE[1][147] ,
         \CACHE[1][146] , \CACHE[1][145] , \CACHE[1][144] , \CACHE[1][143] ,
         \CACHE[1][142] , \CACHE[1][141] , \CACHE[1][140] , \CACHE[1][139] ,
         \CACHE[1][138] , \CACHE[1][137] , \CACHE[1][136] , \CACHE[1][135] ,
         \CACHE[1][134] , \CACHE[1][133] , \CACHE[1][132] , \CACHE[1][131] ,
         \CACHE[1][130] , \CACHE[1][129] , \CACHE[1][128] , \CACHE[1][127] ,
         \CACHE[1][126] , \CACHE[1][125] , \CACHE[1][124] , \CACHE[1][123] ,
         \CACHE[1][122] , \CACHE[1][121] , \CACHE[1][120] , \CACHE[1][119] ,
         \CACHE[1][118] , \CACHE[1][117] , \CACHE[1][116] , \CACHE[1][115] ,
         \CACHE[1][114] , \CACHE[1][113] , \CACHE[1][112] , \CACHE[1][111] ,
         \CACHE[1][110] , \CACHE[1][109] , \CACHE[1][108] , \CACHE[1][107] ,
         \CACHE[1][106] , \CACHE[1][105] , \CACHE[1][104] , \CACHE[1][103] ,
         \CACHE[1][102] , \CACHE[1][101] , \CACHE[1][100] , \CACHE[1][99] ,
         \CACHE[1][98] , \CACHE[1][97] , \CACHE[1][96] , \CACHE[1][95] ,
         \CACHE[1][94] , \CACHE[1][93] , \CACHE[1][92] , \CACHE[1][91] ,
         \CACHE[1][90] , \CACHE[1][89] , \CACHE[1][88] , \CACHE[1][87] ,
         \CACHE[1][86] , \CACHE[1][85] , \CACHE[1][84] , \CACHE[1][83] ,
         \CACHE[1][82] , \CACHE[1][81] , \CACHE[1][80] , \CACHE[1][79] ,
         \CACHE[1][78] , \CACHE[1][77] , \CACHE[1][76] , \CACHE[1][75] ,
         \CACHE[1][74] , \CACHE[1][73] , \CACHE[1][72] , \CACHE[1][71] ,
         \CACHE[1][70] , \CACHE[1][69] , \CACHE[1][68] , \CACHE[1][67] ,
         \CACHE[1][66] , \CACHE[1][65] , \CACHE[1][64] , \CACHE[1][63] ,
         \CACHE[1][62] , \CACHE[1][61] , \CACHE[1][60] , \CACHE[1][59] ,
         \CACHE[1][58] , \CACHE[1][57] , \CACHE[1][56] , \CACHE[1][55] ,
         \CACHE[1][54] , \CACHE[1][53] , \CACHE[1][52] , \CACHE[1][51] ,
         \CACHE[1][50] , \CACHE[1][49] , \CACHE[1][48] , \CACHE[1][47] ,
         \CACHE[1][46] , \CACHE[1][45] , \CACHE[1][44] , \CACHE[1][43] ,
         \CACHE[1][42] , \CACHE[1][41] , \CACHE[1][40] , \CACHE[1][39] ,
         \CACHE[1][38] , \CACHE[1][37] , \CACHE[1][36] , \CACHE[1][35] ,
         \CACHE[1][34] , \CACHE[1][33] , \CACHE[1][32] , \CACHE[1][31] ,
         \CACHE[1][30] , \CACHE[1][29] , \CACHE[1][28] , \CACHE[1][27] ,
         \CACHE[1][26] , \CACHE[1][25] , \CACHE[1][24] , \CACHE[1][23] ,
         \CACHE[1][22] , \CACHE[1][21] , \CACHE[1][20] , \CACHE[1][19] ,
         \CACHE[1][18] , \CACHE[1][17] , \CACHE[1][16] , \CACHE[1][15] ,
         \CACHE[1][14] , \CACHE[1][13] , \CACHE[1][12] , \CACHE[1][11] ,
         \CACHE[1][10] , \CACHE[1][9] , \CACHE[1][8] , \CACHE[1][7] ,
         \CACHE[1][6] , \CACHE[1][5] , \CACHE[1][4] , \CACHE[1][3] ,
         \CACHE[1][2] , \CACHE[1][1] , \CACHE[1][0] , \CACHE[0][154] ,
         \CACHE[0][153] , \CACHE[0][152] , \CACHE[0][151] , \CACHE[0][150] ,
         \CACHE[0][149] , \CACHE[0][148] , \CACHE[0][147] , \CACHE[0][146] ,
         \CACHE[0][145] , \CACHE[0][144] , \CACHE[0][143] , \CACHE[0][142] ,
         \CACHE[0][141] , \CACHE[0][140] , \CACHE[0][139] , \CACHE[0][138] ,
         \CACHE[0][137] , \CACHE[0][136] , \CACHE[0][135] , \CACHE[0][134] ,
         \CACHE[0][133] , \CACHE[0][132] , \CACHE[0][131] , \CACHE[0][130] ,
         \CACHE[0][129] , \CACHE[0][128] , \CACHE[0][127] , \CACHE[0][126] ,
         \CACHE[0][125] , \CACHE[0][124] , \CACHE[0][123] , \CACHE[0][122] ,
         \CACHE[0][121] , \CACHE[0][120] , \CACHE[0][119] , \CACHE[0][118] ,
         \CACHE[0][117] , \CACHE[0][116] , \CACHE[0][115] , \CACHE[0][114] ,
         \CACHE[0][113] , \CACHE[0][112] , \CACHE[0][111] , \CACHE[0][110] ,
         \CACHE[0][109] , \CACHE[0][108] , \CACHE[0][107] , \CACHE[0][106] ,
         \CACHE[0][105] , \CACHE[0][104] , \CACHE[0][103] , \CACHE[0][102] ,
         \CACHE[0][101] , \CACHE[0][100] , \CACHE[0][99] , \CACHE[0][98] ,
         \CACHE[0][97] , \CACHE[0][96] , \CACHE[0][95] , \CACHE[0][94] ,
         \CACHE[0][93] , \CACHE[0][92] , \CACHE[0][91] , \CACHE[0][90] ,
         \CACHE[0][89] , \CACHE[0][88] , \CACHE[0][87] , \CACHE[0][86] ,
         \CACHE[0][85] , \CACHE[0][84] , \CACHE[0][83] , \CACHE[0][82] ,
         \CACHE[0][81] , \CACHE[0][80] , \CACHE[0][79] , \CACHE[0][78] ,
         \CACHE[0][77] , \CACHE[0][76] , \CACHE[0][75] , \CACHE[0][74] ,
         \CACHE[0][73] , \CACHE[0][72] , \CACHE[0][71] , \CACHE[0][70] ,
         \CACHE[0][69] , \CACHE[0][68] , \CACHE[0][67] , \CACHE[0][66] ,
         \CACHE[0][65] , \CACHE[0][64] , \CACHE[0][63] , \CACHE[0][62] ,
         \CACHE[0][61] , \CACHE[0][60] , \CACHE[0][59] , \CACHE[0][58] ,
         \CACHE[0][57] , \CACHE[0][56] , \CACHE[0][55] , \CACHE[0][54] ,
         \CACHE[0][53] , \CACHE[0][52] , \CACHE[0][51] , \CACHE[0][50] ,
         \CACHE[0][49] , \CACHE[0][48] , \CACHE[0][47] , \CACHE[0][46] ,
         \CACHE[0][45] , \CACHE[0][44] , \CACHE[0][43] , \CACHE[0][42] ,
         \CACHE[0][41] , \CACHE[0][40] , \CACHE[0][39] , \CACHE[0][38] ,
         \CACHE[0][37] , \CACHE[0][36] , \CACHE[0][35] , \CACHE[0][34] ,
         \CACHE[0][33] , \CACHE[0][32] , \CACHE[0][31] , \CACHE[0][30] ,
         \CACHE[0][29] , \CACHE[0][28] , \CACHE[0][27] , \CACHE[0][26] ,
         \CACHE[0][25] , \CACHE[0][24] , \CACHE[0][23] , \CACHE[0][22] ,
         \CACHE[0][21] , \CACHE[0][20] , \CACHE[0][19] , \CACHE[0][18] ,
         \CACHE[0][17] , \CACHE[0][16] , \CACHE[0][15] , \CACHE[0][14] ,
         \CACHE[0][13] , \CACHE[0][12] , \CACHE[0][11] , \CACHE[0][10] ,
         \CACHE[0][9] , \CACHE[0][8] , \CACHE[0][7] , \CACHE[0][6] ,
         \CACHE[0][5] , \CACHE[0][4] , \CACHE[0][3] , \CACHE[0][2] ,
         \CACHE[0][1] , \CACHE[0][0] , N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96,
         N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108,
         N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119,
         N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130,
         N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141,
         N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152,
         N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163,
         N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174,
         N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185,
         N186, N187, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n313, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n3020, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280;
  assign N30 = proc_addr[2];
  assign N31 = proc_addr[3];
  assign N32 = proc_addr[4];

  DFFRX1 \CACHE_reg[7][154]  ( .D(n3801), .CK(clk), .RN(n3057), .Q(
        \CACHE[7][154] ), .QN(n5041) );
  DFFRX1 \CACHE_reg[7][153]  ( .D(n3802), .CK(clk), .RN(n3057), .Q(
        \CACHE[7][153] ), .QN(n5042) );
  DFFRX1 \CACHE_reg[7][152]  ( .D(n3803), .CK(clk), .RN(n474), .Q(
        \CACHE[7][152] ), .QN(n5043) );
  DFFRX1 \CACHE_reg[7][151]  ( .D(n3804), .CK(clk), .RN(n475), .Q(
        \CACHE[7][151] ), .QN(n5044) );
  DFFRX1 \CACHE_reg[7][150]  ( .D(n3805), .CK(clk), .RN(n476), .Q(
        \CACHE[7][150] ), .QN(n5045) );
  DFFRX1 \CACHE_reg[7][149]  ( .D(n3806), .CK(clk), .RN(n476), .Q(
        \CACHE[7][149] ), .QN(n5046) );
  DFFRX1 \CACHE_reg[7][148]  ( .D(n3807), .CK(clk), .RN(n477), .Q(
        \CACHE[7][148] ), .QN(n5047) );
  DFFRX1 \CACHE_reg[7][147]  ( .D(n3808), .CK(clk), .RN(n478), .Q(
        \CACHE[7][147] ), .QN(n5048) );
  DFFRX1 \CACHE_reg[7][146]  ( .D(n3809), .CK(clk), .RN(n478), .Q(
        \CACHE[7][146] ), .QN(n5049) );
  DFFRX1 \CACHE_reg[7][145]  ( .D(n3810), .CK(clk), .RN(n479), .Q(
        \CACHE[7][145] ), .QN(n5050) );
  DFFRX1 \CACHE_reg[7][144]  ( .D(n3811), .CK(clk), .RN(n480), .Q(
        \CACHE[7][144] ), .QN(n5051) );
  DFFRX1 \CACHE_reg[7][143]  ( .D(n3812), .CK(clk), .RN(n480), .Q(
        \CACHE[7][143] ), .QN(n5052) );
  DFFRX1 \CACHE_reg[7][142]  ( .D(n3813), .CK(clk), .RN(n481), .Q(
        \CACHE[7][142] ), .QN(n5053) );
  DFFRX1 \CACHE_reg[7][141]  ( .D(n3814), .CK(clk), .RN(n482), .Q(
        \CACHE[7][141] ), .QN(n5054) );
  DFFRX1 \CACHE_reg[7][140]  ( .D(n3815), .CK(clk), .RN(n482), .Q(
        \CACHE[7][140] ), .QN(n5055) );
  DFFRX1 \CACHE_reg[7][139]  ( .D(n3816), .CK(clk), .RN(n490), .Q(
        \CACHE[7][139] ), .QN(n5056) );
  DFFRX1 \CACHE_reg[7][138]  ( .D(n3817), .CK(clk), .RN(n483), .Q(
        \CACHE[7][138] ), .QN(n5057) );
  DFFRX1 \CACHE_reg[7][137]  ( .D(n3818), .CK(clk), .RN(n484), .Q(
        \CACHE[7][137] ), .QN(n5058) );
  DFFRX1 \CACHE_reg[7][136]  ( .D(n3819), .CK(clk), .RN(n484), .Q(
        \CACHE[7][136] ), .QN(n5059) );
  DFFRX1 \CACHE_reg[7][135]  ( .D(n3820), .CK(clk), .RN(n485), .Q(
        \CACHE[7][135] ), .QN(n5060) );
  DFFRX1 \CACHE_reg[7][134]  ( .D(n3821), .CK(clk), .RN(n486), .Q(
        \CACHE[7][134] ), .QN(n5061) );
  DFFRX1 \CACHE_reg[7][133]  ( .D(n3822), .CK(clk), .RN(n486), .Q(
        \CACHE[7][133] ), .QN(n5062) );
  DFFRX1 \CACHE_reg[7][132]  ( .D(n3823), .CK(clk), .RN(n474), .Q(
        \CACHE[7][132] ), .QN(n5063) );
  DFFRX1 \CACHE_reg[7][131]  ( .D(n3824), .CK(clk), .RN(n487), .Q(
        \CACHE[7][131] ), .QN(n5064) );
  DFFRX1 \CACHE_reg[7][130]  ( .D(n3825), .CK(clk), .RN(n488), .Q(
        \CACHE[7][130] ), .QN(n5065) );
  DFFRX1 \CACHE_reg[7][129]  ( .D(n3826), .CK(clk), .RN(n488), .Q(
        \CACHE[7][129] ), .QN(n5066) );
  DFFRX1 \CACHE_reg[7][128]  ( .D(n3827), .CK(clk), .RN(n489), .Q(
        \CACHE[7][128] ), .QN(n5067) );
  DFFRX1 \CACHE_reg[7][127]  ( .D(n3828), .CK(clk), .RN(n3057), .Q(
        \CACHE[7][127] ), .QN(n5068) );
  DFFRX1 \CACHE_reg[7][126]  ( .D(n3829), .CK(clk), .RN(n491), .Q(
        \CACHE[7][126] ), .QN(n5069) );
  DFFRX1 \CACHE_reg[7][125]  ( .D(n3830), .CK(clk), .RN(n533), .Q(
        \CACHE[7][125] ), .QN(n5070) );
  DFFRX1 \CACHE_reg[7][124]  ( .D(n3831), .CK(clk), .RN(n534), .Q(
        \CACHE[7][124] ), .QN(n5071) );
  DFFRX1 \CACHE_reg[7][123]  ( .D(n3832), .CK(clk), .RN(n535), .Q(
        \CACHE[7][123] ), .QN(n5072) );
  DFFRX1 \CACHE_reg[7][122]  ( .D(n3833), .CK(clk), .RN(n535), .Q(
        \CACHE[7][122] ), .QN(n5073) );
  DFFRX1 \CACHE_reg[7][121]  ( .D(n3834), .CK(clk), .RN(n536), .Q(
        \CACHE[7][121] ), .QN(n5074) );
  DFFRX1 \CACHE_reg[7][120]  ( .D(n3835), .CK(clk), .RN(n537), .Q(
        \CACHE[7][120] ), .QN(n5075) );
  DFFRX1 \CACHE_reg[7][119]  ( .D(n3836), .CK(clk), .RN(n537), .Q(
        \CACHE[7][119] ), .QN(n5076) );
  DFFRX1 \CACHE_reg[7][118]  ( .D(n3837), .CK(clk), .RN(n538), .Q(
        \CACHE[7][118] ), .QN(n5077) );
  DFFRX1 \CACHE_reg[7][117]  ( .D(n3838), .CK(clk), .RN(n539), .Q(
        \CACHE[7][117] ), .QN(n5078) );
  DFFRX1 \CACHE_reg[7][116]  ( .D(n3839), .CK(clk), .RN(n539), .Q(
        \CACHE[7][116] ), .QN(n5079) );
  DFFRX1 \CACHE_reg[7][115]  ( .D(n3840), .CK(clk), .RN(n540), .Q(
        \CACHE[7][115] ), .QN(n5080) );
  DFFRX1 \CACHE_reg[7][114]  ( .D(n3841), .CK(clk), .RN(n3020), .Q(
        \CACHE[7][114] ), .QN(n5081) );
  DFFRX1 \CACHE_reg[7][113]  ( .D(n3842), .CK(clk), .RN(n3020), .Q(
        \CACHE[7][113] ), .QN(n5082) );
  DFFRX1 \CACHE_reg[7][112]  ( .D(n3843), .CK(clk), .RN(n3022), .Q(
        \CACHE[7][112] ), .QN(n5083) );
  DFFRX1 \CACHE_reg[7][111]  ( .D(n3844), .CK(clk), .RN(n3023), .Q(
        \CACHE[7][111] ), .QN(n5084) );
  DFFRX1 \CACHE_reg[7][110]  ( .D(n3845), .CK(clk), .RN(n3023), .Q(
        \CACHE[7][110] ), .QN(n5085) );
  DFFRX1 \CACHE_reg[7][109]  ( .D(n3846), .CK(clk), .RN(n3024), .Q(
        \CACHE[7][109] ), .QN(n5086) );
  DFFRX1 \CACHE_reg[7][108]  ( .D(n3847), .CK(clk), .RN(n3025), .Q(
        \CACHE[7][108] ), .QN(n5087) );
  DFFRX1 \CACHE_reg[7][107]  ( .D(n3848), .CK(clk), .RN(n3025), .Q(
        \CACHE[7][107] ), .QN(n5088) );
  DFFRX1 \CACHE_reg[7][106]  ( .D(n3849), .CK(clk), .RN(n3026), .Q(
        \CACHE[7][106] ), .QN(n5089) );
  DFFRX1 \CACHE_reg[7][105]  ( .D(n3850), .CK(clk), .RN(n3027), .Q(
        \CACHE[7][105] ), .QN(n5090) );
  DFFRX1 \CACHE_reg[7][104]  ( .D(n3851), .CK(clk), .RN(n3027), .Q(
        \CACHE[7][104] ), .QN(n5091) );
  DFFRX1 \CACHE_reg[7][103]  ( .D(n3852), .CK(clk), .RN(n3028), .Q(
        \CACHE[7][103] ), .QN(n5092) );
  DFFRX1 \CACHE_reg[7][102]  ( .D(n3853), .CK(clk), .RN(n3029), .Q(
        \CACHE[7][102] ), .QN(n5093) );
  DFFRX1 \CACHE_reg[7][101]  ( .D(n3854), .CK(clk), .RN(n3029), .Q(
        \CACHE[7][101] ), .QN(n5094) );
  DFFRX1 \CACHE_reg[7][100]  ( .D(n3855), .CK(clk), .RN(n3030), .Q(
        \CACHE[7][100] ), .QN(n5095) );
  DFFRX1 \CACHE_reg[7][99]  ( .D(n3856), .CK(clk), .RN(n3031), .Q(
        \CACHE[7][99] ), .QN(n5096) );
  DFFRX1 \CACHE_reg[7][98]  ( .D(n3857), .CK(clk), .RN(n3031), .Q(
        \CACHE[7][98] ), .QN(n5097) );
  DFFRX1 \CACHE_reg[7][97]  ( .D(n3858), .CK(clk), .RN(n3032), .Q(
        \CACHE[7][97] ), .QN(n5098) );
  DFFRX1 \CACHE_reg[7][96]  ( .D(n3859), .CK(clk), .RN(n3033), .Q(
        \CACHE[7][96] ), .QN(n5099) );
  DFFRX1 \CACHE_reg[7][95]  ( .D(n3860), .CK(clk), .RN(n3033), .Q(
        \CACHE[7][95] ), .QN(n5100) );
  DFFRX1 \CACHE_reg[7][94]  ( .D(n3861), .CK(clk), .RN(n3034), .Q(
        \CACHE[7][94] ), .QN(n5101) );
  DFFRX1 \CACHE_reg[7][93]  ( .D(n3862), .CK(clk), .RN(n3035), .Q(
        \CACHE[7][93] ), .QN(n5102) );
  DFFRX1 \CACHE_reg[7][92]  ( .D(n3863), .CK(clk), .RN(n3035), .Q(
        \CACHE[7][92] ), .QN(n5103) );
  DFFRX1 \CACHE_reg[7][91]  ( .D(n3864), .CK(clk), .RN(n3036), .Q(
        \CACHE[7][91] ), .QN(n5104) );
  DFFRX1 \CACHE_reg[7][90]  ( .D(n3865), .CK(clk), .RN(n3037), .Q(
        \CACHE[7][90] ), .QN(n5105) );
  DFFRX1 \CACHE_reg[7][89]  ( .D(n3866), .CK(clk), .RN(n3037), .Q(
        \CACHE[7][89] ), .QN(n5106) );
  DFFRX1 \CACHE_reg[7][88]  ( .D(n3867), .CK(clk), .RN(n3038), .Q(
        \CACHE[7][88] ), .QN(n5107) );
  DFFRX1 \CACHE_reg[7][87]  ( .D(n3868), .CK(clk), .RN(n3039), .Q(
        \CACHE[7][87] ), .QN(n5108) );
  DFFRX1 \CACHE_reg[7][86]  ( .D(n3869), .CK(clk), .RN(n3039), .Q(
        \CACHE[7][86] ), .QN(n5109) );
  DFFRX1 \CACHE_reg[7][85]  ( .D(n3870), .CK(clk), .RN(n3040), .Q(
        \CACHE[7][85] ), .QN(n5110) );
  DFFRX1 \CACHE_reg[7][84]  ( .D(n3871), .CK(clk), .RN(n3041), .Q(
        \CACHE[7][84] ), .QN(n5111) );
  DFFRX1 \CACHE_reg[7][83]  ( .D(n3872), .CK(clk), .RN(n3041), .Q(
        \CACHE[7][83] ), .QN(n5112) );
  DFFRX1 \CACHE_reg[7][82]  ( .D(n3873), .CK(clk), .RN(n3042), .Q(
        \CACHE[7][82] ), .QN(n5113) );
  DFFRX1 \CACHE_reg[7][81]  ( .D(n3874), .CK(clk), .RN(n3043), .Q(
        \CACHE[7][81] ), .QN(n5114) );
  DFFRX1 \CACHE_reg[7][80]  ( .D(n3875), .CK(clk), .RN(n3043), .Q(
        \CACHE[7][80] ), .QN(n5115) );
  DFFRX1 \CACHE_reg[7][79]  ( .D(n3876), .CK(clk), .RN(n3044), .Q(
        \CACHE[7][79] ), .QN(n5116) );
  DFFRX1 \CACHE_reg[7][78]  ( .D(n3877), .CK(clk), .RN(n3045), .Q(
        \CACHE[7][78] ), .QN(n5117) );
  DFFRX1 \CACHE_reg[7][77]  ( .D(n3878), .CK(clk), .RN(n3045), .Q(
        \CACHE[7][77] ), .QN(n5118) );
  DFFRX1 \CACHE_reg[7][76]  ( .D(n3879), .CK(clk), .RN(n3046), .Q(
        \CACHE[7][76] ), .QN(n5119) );
  DFFRX1 \CACHE_reg[7][75]  ( .D(n3880), .CK(clk), .RN(n3047), .Q(
        \CACHE[7][75] ), .QN(n5120) );
  DFFRX1 \CACHE_reg[7][74]  ( .D(n3881), .CK(clk), .RN(n3047), .Q(
        \CACHE[7][74] ), .QN(n5121) );
  DFFRX1 \CACHE_reg[7][73]  ( .D(n3882), .CK(clk), .RN(n3048), .Q(
        \CACHE[7][73] ), .QN(n5122) );
  DFFRX1 \CACHE_reg[7][72]  ( .D(n3883), .CK(clk), .RN(n3049), .Q(
        \CACHE[7][72] ), .QN(n5123) );
  DFFRX1 \CACHE_reg[7][71]  ( .D(n3884), .CK(clk), .RN(n3049), .Q(
        \CACHE[7][71] ), .QN(n5124) );
  DFFRX1 \CACHE_reg[7][70]  ( .D(n3885), .CK(clk), .RN(n3050), .Q(
        \CACHE[7][70] ), .QN(n5125) );
  DFFRX1 \CACHE_reg[7][69]  ( .D(n3886), .CK(clk), .RN(n3051), .Q(
        \CACHE[7][69] ), .QN(n5126) );
  DFFRX1 \CACHE_reg[7][68]  ( .D(n3887), .CK(clk), .RN(n3051), .Q(
        \CACHE[7][68] ), .QN(n5127) );
  DFFRX1 \CACHE_reg[7][67]  ( .D(n3888), .CK(clk), .RN(n3052), .Q(
        \CACHE[7][67] ), .QN(n5128) );
  DFFRX1 \CACHE_reg[7][66]  ( .D(n3889), .CK(clk), .RN(n3053), .Q(
        \CACHE[7][66] ), .QN(n5129) );
  DFFRX1 \CACHE_reg[7][65]  ( .D(n3890), .CK(clk), .RN(n3053), .Q(
        \CACHE[7][65] ), .QN(n5130) );
  DFFRX1 \CACHE_reg[7][64]  ( .D(n3891), .CK(clk), .RN(n3054), .Q(
        \CACHE[7][64] ), .QN(n5131) );
  DFFRX1 \CACHE_reg[7][63]  ( .D(n3892), .CK(clk), .RN(n512), .Q(
        \CACHE[7][63] ), .QN(n5132) );
  DFFRX1 \CACHE_reg[7][62]  ( .D(n3893), .CK(clk), .RN(n513), .Q(
        \CACHE[7][62] ), .QN(n5133) );
  DFFRX1 \CACHE_reg[7][61]  ( .D(n3894), .CK(clk), .RN(n513), .Q(
        \CACHE[7][61] ), .QN(n5134) );
  DFFRX1 \CACHE_reg[7][60]  ( .D(n3895), .CK(clk), .RN(n514), .Q(
        \CACHE[7][60] ), .QN(n5135) );
  DFFRX1 \CACHE_reg[7][59]  ( .D(n3896), .CK(clk), .RN(n515), .Q(
        \CACHE[7][59] ), .QN(n5136) );
  DFFRX1 \CACHE_reg[7][58]  ( .D(n3897), .CK(clk), .RN(n515), .Q(
        \CACHE[7][58] ), .QN(n5137) );
  DFFRX1 \CACHE_reg[7][57]  ( .D(n3898), .CK(clk), .RN(n516), .Q(
        \CACHE[7][57] ), .QN(n5138) );
  DFFRX1 \CACHE_reg[7][56]  ( .D(n3899), .CK(clk), .RN(n517), .Q(
        \CACHE[7][56] ), .QN(n5139) );
  DFFRX1 \CACHE_reg[7][55]  ( .D(n3900), .CK(clk), .RN(n517), .Q(
        \CACHE[7][55] ), .QN(n5140) );
  DFFRX1 \CACHE_reg[7][54]  ( .D(n3901), .CK(clk), .RN(n518), .Q(
        \CACHE[7][54] ), .QN(n5141) );
  DFFRX1 \CACHE_reg[7][53]  ( .D(n3902), .CK(clk), .RN(n519), .Q(
        \CACHE[7][53] ), .QN(n5142) );
  DFFRX1 \CACHE_reg[7][52]  ( .D(n3903), .CK(clk), .RN(n519), .Q(
        \CACHE[7][52] ), .QN(n5143) );
  DFFRX1 \CACHE_reg[7][51]  ( .D(n3904), .CK(clk), .RN(n520), .Q(
        \CACHE[7][51] ), .QN(n5144) );
  DFFRX1 \CACHE_reg[7][50]  ( .D(n3905), .CK(clk), .RN(n521), .Q(
        \CACHE[7][50] ), .QN(n5145) );
  DFFRX1 \CACHE_reg[7][49]  ( .D(n3906), .CK(clk), .RN(n521), .Q(
        \CACHE[7][49] ), .QN(n5146) );
  DFFRX1 \CACHE_reg[7][48]  ( .D(n3907), .CK(clk), .RN(n522), .Q(
        \CACHE[7][48] ), .QN(n5147) );
  DFFRX1 \CACHE_reg[7][47]  ( .D(n3908), .CK(clk), .RN(n523), .Q(
        \CACHE[7][47] ), .QN(n5148) );
  DFFRX1 \CACHE_reg[7][46]  ( .D(n3909), .CK(clk), .RN(n523), .Q(
        \CACHE[7][46] ), .QN(n5149) );
  DFFRX1 \CACHE_reg[7][45]  ( .D(n3910), .CK(clk), .RN(n524), .Q(
        \CACHE[7][45] ), .QN(n5150) );
  DFFRX1 \CACHE_reg[7][44]  ( .D(n3911), .CK(clk), .RN(n525), .Q(
        \CACHE[7][44] ), .QN(n5151) );
  DFFRX1 \CACHE_reg[7][43]  ( .D(n3912), .CK(clk), .RN(n525), .Q(
        \CACHE[7][43] ), .QN(n5152) );
  DFFRX1 \CACHE_reg[7][42]  ( .D(n3913), .CK(clk), .RN(n526), .Q(
        \CACHE[7][42] ), .QN(n5153) );
  DFFRX1 \CACHE_reg[7][41]  ( .D(n3914), .CK(clk), .RN(n527), .Q(
        \CACHE[7][41] ), .QN(n5154) );
  DFFRX1 \CACHE_reg[7][40]  ( .D(n3915), .CK(clk), .RN(n527), .Q(
        \CACHE[7][40] ), .QN(n5155) );
  DFFRX1 \CACHE_reg[7][39]  ( .D(n3916), .CK(clk), .RN(n528), .Q(
        \CACHE[7][39] ), .QN(n5156) );
  DFFRX1 \CACHE_reg[7][38]  ( .D(n3917), .CK(clk), .RN(n529), .Q(
        \CACHE[7][38] ), .QN(n5157) );
  DFFRX1 \CACHE_reg[7][37]  ( .D(n3918), .CK(clk), .RN(n529), .Q(
        \CACHE[7][37] ), .QN(n5158) );
  DFFRX1 \CACHE_reg[7][36]  ( .D(n3919), .CK(clk), .RN(n530), .Q(
        \CACHE[7][36] ), .QN(n5159) );
  DFFRX1 \CACHE_reg[7][35]  ( .D(n3920), .CK(clk), .RN(n531), .Q(
        \CACHE[7][35] ), .QN(n5160) );
  DFFRX1 \CACHE_reg[7][34]  ( .D(n3921), .CK(clk), .RN(n531), .Q(
        \CACHE[7][34] ), .QN(n5161) );
  DFFRX1 \CACHE_reg[7][33]  ( .D(n3922), .CK(clk), .RN(n532), .Q(
        \CACHE[7][33] ), .QN(n5162) );
  DFFRX1 \CACHE_reg[7][32]  ( .D(n3923), .CK(clk), .RN(n533), .Q(
        \CACHE[7][32] ), .QN(n5163) );
  DFFRX1 \CACHE_reg[7][31]  ( .D(n3924), .CK(clk), .RN(n490), .Q(
        \CACHE[7][31] ), .QN(n5164) );
  DFFRX1 \CACHE_reg[7][30]  ( .D(n3925), .CK(clk), .RN(n3057), .Q(
        \CACHE[7][30] ), .QN(n5165) );
  DFFRX1 \CACHE_reg[7][29]  ( .D(n3926), .CK(clk), .RN(n492), .Q(
        \CACHE[7][29] ), .QN(n5166) );
  DFFRX1 \CACHE_reg[7][28]  ( .D(n3927), .CK(clk), .RN(n493), .Q(
        \CACHE[7][28] ), .QN(n5167) );
  DFFRX1 \CACHE_reg[7][27]  ( .D(n3928), .CK(clk), .RN(n493), .Q(
        \CACHE[7][27] ), .QN(n5168) );
  DFFRX1 \CACHE_reg[7][26]  ( .D(n3929), .CK(clk), .RN(n494), .Q(
        \CACHE[7][26] ), .QN(n5169) );
  DFFRX1 \CACHE_reg[7][25]  ( .D(n3930), .CK(clk), .RN(n495), .Q(
        \CACHE[7][25] ), .QN(n5170) );
  DFFRX1 \CACHE_reg[7][24]  ( .D(n3931), .CK(clk), .RN(n495), .Q(
        \CACHE[7][24] ), .QN(n5171) );
  DFFRX1 \CACHE_reg[7][23]  ( .D(n3932), .CK(clk), .RN(n496), .Q(
        \CACHE[7][23] ), .QN(n5172) );
  DFFRX1 \CACHE_reg[7][22]  ( .D(n3933), .CK(clk), .RN(n497), .Q(
        \CACHE[7][22] ), .QN(n5173) );
  DFFRX1 \CACHE_reg[7][21]  ( .D(n3934), .CK(clk), .RN(n497), .Q(
        \CACHE[7][21] ), .QN(n5174) );
  DFFRX1 \CACHE_reg[7][20]  ( .D(n3935), .CK(clk), .RN(n498), .Q(
        \CACHE[7][20] ), .QN(n5175) );
  DFFRX1 \CACHE_reg[7][19]  ( .D(n3936), .CK(clk), .RN(n499), .Q(
        \CACHE[7][19] ), .QN(n5176) );
  DFFRX1 \CACHE_reg[7][18]  ( .D(n3937), .CK(clk), .RN(n499), .Q(
        \CACHE[7][18] ), .QN(n5177) );
  DFFRX1 \CACHE_reg[7][17]  ( .D(n3938), .CK(clk), .RN(n500), .Q(
        \CACHE[7][17] ), .QN(n5178) );
  DFFRX1 \CACHE_reg[7][16]  ( .D(n3939), .CK(clk), .RN(n501), .Q(
        \CACHE[7][16] ), .QN(n5179) );
  DFFRX1 \CACHE_reg[7][15]  ( .D(n3940), .CK(clk), .RN(n501), .Q(
        \CACHE[7][15] ), .QN(n5180) );
  DFFRX1 \CACHE_reg[7][14]  ( .D(n3941), .CK(clk), .RN(n502), .Q(
        \CACHE[7][14] ), .QN(n5181) );
  DFFRX1 \CACHE_reg[7][13]  ( .D(n3942), .CK(clk), .RN(n503), .Q(
        \CACHE[7][13] ), .QN(n5182) );
  DFFRX1 \CACHE_reg[7][12]  ( .D(n3943), .CK(clk), .RN(n503), .Q(
        \CACHE[7][12] ), .QN(n5183) );
  DFFRX1 \CACHE_reg[7][11]  ( .D(n3944), .CK(clk), .RN(n504), .Q(
        \CACHE[7][11] ), .QN(n5184) );
  DFFRX1 \CACHE_reg[7][10]  ( .D(n3945), .CK(clk), .RN(n505), .Q(
        \CACHE[7][10] ), .QN(n5185) );
  DFFRX1 \CACHE_reg[7][9]  ( .D(n3946), .CK(clk), .RN(n505), .Q(\CACHE[7][9] ), 
        .QN(n5186) );
  DFFRX1 \CACHE_reg[7][8]  ( .D(n3947), .CK(clk), .RN(n506), .Q(\CACHE[7][8] ), 
        .QN(n5187) );
  DFFRX1 \CACHE_reg[7][7]  ( .D(n3948), .CK(clk), .RN(n507), .Q(\CACHE[7][7] ), 
        .QN(n5188) );
  DFFRX1 \CACHE_reg[7][6]  ( .D(n3949), .CK(clk), .RN(n507), .Q(\CACHE[7][6] ), 
        .QN(n5189) );
  DFFRX1 \CACHE_reg[7][5]  ( .D(n3950), .CK(clk), .RN(n508), .Q(\CACHE[7][5] ), 
        .QN(n5190) );
  DFFRX1 \CACHE_reg[7][4]  ( .D(n3951), .CK(clk), .RN(n509), .Q(\CACHE[7][4] ), 
        .QN(n5191) );
  DFFRX1 \CACHE_reg[7][3]  ( .D(n3952), .CK(clk), .RN(n509), .Q(\CACHE[7][3] ), 
        .QN(n5192) );
  DFFRX1 \CACHE_reg[7][2]  ( .D(n3953), .CK(clk), .RN(n510), .Q(\CACHE[7][2] ), 
        .QN(n5193) );
  DFFRX1 \CACHE_reg[7][1]  ( .D(n3954), .CK(clk), .RN(n511), .Q(\CACHE[7][1] ), 
        .QN(n5194) );
  DFFRX1 \CACHE_reg[7][0]  ( .D(n3955), .CK(clk), .RN(n511), .Q(\CACHE[7][0] ), 
        .QN(n5195) );
  DFFRX1 \CACHE_reg[3][154]  ( .D(n4421), .CK(clk), .RN(n3055), .Q(
        \CACHE[3][154] ), .QN(n5661) );
  DFFRX1 \CACHE_reg[3][153]  ( .D(n4422), .CK(clk), .RN(n3055), .Q(
        \CACHE[3][153] ), .QN(n5662) );
  DFFRX1 \CACHE_reg[3][152]  ( .D(n4423), .CK(clk), .RN(n475), .Q(
        \CACHE[3][152] ), .QN(n5663) );
  DFFRX1 \CACHE_reg[3][151]  ( .D(n4424), .CK(clk), .RN(n475), .Q(
        \CACHE[3][151] ), .QN(n5664) );
  DFFRX1 \CACHE_reg[3][150]  ( .D(n4425), .CK(clk), .RN(n476), .Q(
        \CACHE[3][150] ), .QN(n5665) );
  DFFRX1 \CACHE_reg[3][149]  ( .D(n4426), .CK(clk), .RN(n477), .Q(
        \CACHE[3][149] ), .QN(n5666) );
  DFFRX1 \CACHE_reg[3][148]  ( .D(n4427), .CK(clk), .RN(n477), .Q(
        \CACHE[3][148] ), .QN(n5667) );
  DFFRX1 \CACHE_reg[3][147]  ( .D(n4428), .CK(clk), .RN(n478), .Q(
        \CACHE[3][147] ), .QN(n5668) );
  DFFRX1 \CACHE_reg[3][146]  ( .D(n4429), .CK(clk), .RN(n479), .Q(
        \CACHE[3][146] ), .QN(n5669) );
  DFFRX1 \CACHE_reg[3][145]  ( .D(n4430), .CK(clk), .RN(n479), .Q(
        \CACHE[3][145] ), .QN(n5670) );
  DFFRX1 \CACHE_reg[3][144]  ( .D(n4431), .CK(clk), .RN(n480), .Q(
        \CACHE[3][144] ), .QN(n5671) );
  DFFRX1 \CACHE_reg[3][143]  ( .D(n4432), .CK(clk), .RN(n481), .Q(
        \CACHE[3][143] ), .QN(n5672) );
  DFFRX1 \CACHE_reg[3][142]  ( .D(n4433), .CK(clk), .RN(n481), .Q(
        \CACHE[3][142] ), .QN(n5673) );
  DFFRX1 \CACHE_reg[3][141]  ( .D(n4434), .CK(clk), .RN(n482), .Q(
        \CACHE[3][141] ), .QN(n5674) );
  DFFRX1 \CACHE_reg[3][140]  ( .D(n4435), .CK(clk), .RN(n483), .Q(
        \CACHE[3][140] ), .QN(n5675) );
  DFFRX1 \CACHE_reg[3][139]  ( .D(n4436), .CK(clk), .RN(n490), .Q(
        \CACHE[3][139] ), .QN(n5676) );
  DFFRX1 \CACHE_reg[3][138]  ( .D(n4437), .CK(clk), .RN(n483), .Q(
        \CACHE[3][138] ), .QN(n5677) );
  DFFRX1 \CACHE_reg[3][137]  ( .D(n4438), .CK(clk), .RN(n484), .Q(
        \CACHE[3][137] ), .QN(n5678) );
  DFFRX1 \CACHE_reg[3][136]  ( .D(n4439), .CK(clk), .RN(n485), .Q(
        \CACHE[3][136] ), .QN(n5679) );
  DFFRX1 \CACHE_reg[3][135]  ( .D(n4440), .CK(clk), .RN(n485), .Q(
        \CACHE[3][135] ), .QN(n5680) );
  DFFRX1 \CACHE_reg[3][134]  ( .D(n4441), .CK(clk), .RN(n486), .Q(
        \CACHE[3][134] ), .QN(n5681) );
  DFFRX1 \CACHE_reg[3][133]  ( .D(n4442), .CK(clk), .RN(n487), .Q(
        \CACHE[3][133] ), .QN(n5682) );
  DFFRX1 \CACHE_reg[3][132]  ( .D(n4443), .CK(clk), .RN(n474), .Q(
        \CACHE[3][132] ), .QN(n5683) );
  DFFRX1 \CACHE_reg[3][131]  ( .D(n4444), .CK(clk), .RN(n487), .Q(
        \CACHE[3][131] ), .QN(n5684) );
  DFFRX1 \CACHE_reg[3][130]  ( .D(n4445), .CK(clk), .RN(n488), .Q(
        \CACHE[3][130] ), .QN(n5685) );
  DFFRX1 \CACHE_reg[3][129]  ( .D(n4446), .CK(clk), .RN(n489), .Q(
        \CACHE[3][129] ), .QN(n5686) );
  DFFRX1 \CACHE_reg[3][128]  ( .D(n4447), .CK(clk), .RN(n489), .Q(
        \CACHE[3][128] ), .QN(n5687) );
  DFFRX1 \CACHE_reg[3][127]  ( .D(n4448), .CK(clk), .RN(n3055), .Q(
        \CACHE[3][127] ), .QN(n5688) );
  DFFRX1 \CACHE_reg[3][126]  ( .D(n4449), .CK(clk), .RN(n491), .Q(
        \CACHE[3][126] ), .QN(n5689) );
  DFFRX1 \CACHE_reg[3][125]  ( .D(n4450), .CK(clk), .RN(n534), .Q(
        \CACHE[3][125] ), .QN(n5690) );
  DFFRX1 \CACHE_reg[3][124]  ( .D(n4451), .CK(clk), .RN(n534), .Q(
        \CACHE[3][124] ), .QN(n5691) );
  DFFRX1 \CACHE_reg[3][123]  ( .D(n4452), .CK(clk), .RN(n535), .Q(
        \CACHE[3][123] ), .QN(n5692) );
  DFFRX1 \CACHE_reg[3][122]  ( .D(n4453), .CK(clk), .RN(n536), .Q(
        \CACHE[3][122] ), .QN(n5693) );
  DFFRX1 \CACHE_reg[3][121]  ( .D(n4454), .CK(clk), .RN(n536), .Q(
        \CACHE[3][121] ), .QN(n5694) );
  DFFRX1 \CACHE_reg[3][120]  ( .D(n4455), .CK(clk), .RN(n537), .Q(
        \CACHE[3][120] ), .QN(n5695) );
  DFFRX1 \CACHE_reg[3][119]  ( .D(n4456), .CK(clk), .RN(n538), .Q(
        \CACHE[3][119] ), .QN(n5696) );
  DFFRX1 \CACHE_reg[3][118]  ( .D(n4457), .CK(clk), .RN(n538), .Q(
        \CACHE[3][118] ), .QN(n5697) );
  DFFRX1 \CACHE_reg[3][117]  ( .D(n4458), .CK(clk), .RN(n539), .Q(
        \CACHE[3][117] ), .QN(n5698) );
  DFFRX1 \CACHE_reg[3][116]  ( .D(n4459), .CK(clk), .RN(n540), .Q(
        \CACHE[3][116] ), .QN(n5699) );
  DFFRX1 \CACHE_reg[3][115]  ( .D(n4460), .CK(clk), .RN(n540), .Q(
        \CACHE[3][115] ), .QN(n5700) );
  DFFRX1 \CACHE_reg[3][114]  ( .D(n4461), .CK(clk), .RN(n3020), .Q(
        \CACHE[3][114] ), .QN(n5701) );
  DFFRX1 \CACHE_reg[3][113]  ( .D(n4462), .CK(clk), .RN(n3022), .Q(
        \CACHE[3][113] ), .QN(n5702) );
  DFFRX1 \CACHE_reg[3][112]  ( .D(n4463), .CK(clk), .RN(n3022), .Q(
        \CACHE[3][112] ), .QN(n5703) );
  DFFRX1 \CACHE_reg[3][111]  ( .D(n4464), .CK(clk), .RN(n3023), .Q(
        \CACHE[3][111] ), .QN(n5704) );
  DFFRX1 \CACHE_reg[3][110]  ( .D(n4465), .CK(clk), .RN(n3024), .Q(
        \CACHE[3][110] ), .QN(n5705) );
  DFFRX1 \CACHE_reg[3][109]  ( .D(n4466), .CK(clk), .RN(n3024), .Q(
        \CACHE[3][109] ), .QN(n5706) );
  DFFRX1 \CACHE_reg[3][108]  ( .D(n4467), .CK(clk), .RN(n3025), .Q(
        \CACHE[3][108] ), .QN(n5707) );
  DFFRX1 \CACHE_reg[3][107]  ( .D(n4468), .CK(clk), .RN(n3026), .Q(
        \CACHE[3][107] ), .QN(n5708) );
  DFFRX1 \CACHE_reg[3][106]  ( .D(n4469), .CK(clk), .RN(n3026), .Q(
        \CACHE[3][106] ), .QN(n5709) );
  DFFRX1 \CACHE_reg[3][105]  ( .D(n4470), .CK(clk), .RN(n3027), .Q(
        \CACHE[3][105] ), .QN(n5710) );
  DFFRX1 \CACHE_reg[3][104]  ( .D(n4471), .CK(clk), .RN(n3028), .Q(
        \CACHE[3][104] ), .QN(n5711) );
  DFFRX1 \CACHE_reg[3][103]  ( .D(n4472), .CK(clk), .RN(n3028), .Q(
        \CACHE[3][103] ), .QN(n5712) );
  DFFRX1 \CACHE_reg[3][102]  ( .D(n4473), .CK(clk), .RN(n3029), .Q(
        \CACHE[3][102] ), .QN(n5713) );
  DFFRX1 \CACHE_reg[3][101]  ( .D(n4474), .CK(clk), .RN(n3030), .Q(
        \CACHE[3][101] ), .QN(n5714) );
  DFFRX1 \CACHE_reg[3][100]  ( .D(n4475), .CK(clk), .RN(n3030), .Q(
        \CACHE[3][100] ), .QN(n5715) );
  DFFRX1 \CACHE_reg[3][99]  ( .D(n4476), .CK(clk), .RN(n3031), .Q(
        \CACHE[3][99] ), .QN(n5716) );
  DFFRX1 \CACHE_reg[3][98]  ( .D(n4477), .CK(clk), .RN(n3032), .Q(
        \CACHE[3][98] ), .QN(n5717) );
  DFFRX1 \CACHE_reg[3][97]  ( .D(n4478), .CK(clk), .RN(n3032), .Q(
        \CACHE[3][97] ), .QN(n5718) );
  DFFRX1 \CACHE_reg[3][96]  ( .D(n4479), .CK(clk), .RN(n3033), .Q(
        \CACHE[3][96] ), .QN(n5719) );
  DFFRX1 \CACHE_reg[3][95]  ( .D(n4480), .CK(clk), .RN(n3034), .Q(
        \CACHE[3][95] ), .QN(n5720) );
  DFFRX1 \CACHE_reg[3][94]  ( .D(n4481), .CK(clk), .RN(n3034), .Q(
        \CACHE[3][94] ), .QN(n5721) );
  DFFRX1 \CACHE_reg[3][93]  ( .D(n4482), .CK(clk), .RN(n3035), .Q(
        \CACHE[3][93] ), .QN(n5722) );
  DFFRX1 \CACHE_reg[3][92]  ( .D(n4483), .CK(clk), .RN(n3036), .Q(
        \CACHE[3][92] ), .QN(n5723) );
  DFFRX1 \CACHE_reg[3][91]  ( .D(n4484), .CK(clk), .RN(n3036), .Q(
        \CACHE[3][91] ), .QN(n5724) );
  DFFRX1 \CACHE_reg[3][90]  ( .D(n4485), .CK(clk), .RN(n3037), .Q(
        \CACHE[3][90] ), .QN(n5725) );
  DFFRX1 \CACHE_reg[3][89]  ( .D(n4486), .CK(clk), .RN(n3038), .Q(
        \CACHE[3][89] ), .QN(n5726) );
  DFFRX1 \CACHE_reg[3][88]  ( .D(n4487), .CK(clk), .RN(n3038), .Q(
        \CACHE[3][88] ), .QN(n5727) );
  DFFRX1 \CACHE_reg[3][87]  ( .D(n4488), .CK(clk), .RN(n3039), .Q(
        \CACHE[3][87] ), .QN(n5728) );
  DFFRX1 \CACHE_reg[3][86]  ( .D(n4489), .CK(clk), .RN(n3040), .Q(
        \CACHE[3][86] ), .QN(n5729) );
  DFFRX1 \CACHE_reg[3][85]  ( .D(n4490), .CK(clk), .RN(n3040), .Q(
        \CACHE[3][85] ), .QN(n5730) );
  DFFRX1 \CACHE_reg[3][84]  ( .D(n4491), .CK(clk), .RN(n3041), .Q(
        \CACHE[3][84] ), .QN(n5731) );
  DFFRX1 \CACHE_reg[3][83]  ( .D(n4492), .CK(clk), .RN(n3042), .Q(
        \CACHE[3][83] ), .QN(n5732) );
  DFFRX1 \CACHE_reg[3][82]  ( .D(n4493), .CK(clk), .RN(n3042), .Q(
        \CACHE[3][82] ), .QN(n5733) );
  DFFRX1 \CACHE_reg[3][81]  ( .D(n4494), .CK(clk), .RN(n3043), .Q(
        \CACHE[3][81] ), .QN(n5734) );
  DFFRX1 \CACHE_reg[3][80]  ( .D(n4495), .CK(clk), .RN(n3044), .Q(
        \CACHE[3][80] ), .QN(n5735) );
  DFFRX1 \CACHE_reg[3][79]  ( .D(n4496), .CK(clk), .RN(n3044), .Q(
        \CACHE[3][79] ), .QN(n5736) );
  DFFRX1 \CACHE_reg[3][78]  ( .D(n4497), .CK(clk), .RN(n3045), .Q(
        \CACHE[3][78] ), .QN(n5737) );
  DFFRX1 \CACHE_reg[3][77]  ( .D(n4498), .CK(clk), .RN(n3046), .Q(
        \CACHE[3][77] ), .QN(n5738) );
  DFFRX1 \CACHE_reg[3][76]  ( .D(n4499), .CK(clk), .RN(n3046), .Q(
        \CACHE[3][76] ), .QN(n5739) );
  DFFRX1 \CACHE_reg[3][75]  ( .D(n4500), .CK(clk), .RN(n3047), .Q(
        \CACHE[3][75] ), .QN(n5740) );
  DFFRX1 \CACHE_reg[3][74]  ( .D(n4501), .CK(clk), .RN(n3048), .Q(
        \CACHE[3][74] ), .QN(n5741) );
  DFFRX1 \CACHE_reg[3][73]  ( .D(n4502), .CK(clk), .RN(n3048), .Q(
        \CACHE[3][73] ), .QN(n5742) );
  DFFRX1 \CACHE_reg[3][72]  ( .D(n4503), .CK(clk), .RN(n3049), .Q(
        \CACHE[3][72] ), .QN(n5743) );
  DFFRX1 \CACHE_reg[3][71]  ( .D(n4504), .CK(clk), .RN(n3050), .Q(
        \CACHE[3][71] ), .QN(n5744) );
  DFFRX1 \CACHE_reg[3][70]  ( .D(n4505), .CK(clk), .RN(n3050), .Q(
        \CACHE[3][70] ), .QN(n5745) );
  DFFRX1 \CACHE_reg[3][69]  ( .D(n4506), .CK(clk), .RN(n3051), .Q(
        \CACHE[3][69] ), .QN(n5746) );
  DFFRX1 \CACHE_reg[3][68]  ( .D(n4507), .CK(clk), .RN(n3052), .Q(
        \CACHE[3][68] ), .QN(n5747) );
  DFFRX1 \CACHE_reg[3][67]  ( .D(n4508), .CK(clk), .RN(n3052), .Q(
        \CACHE[3][67] ), .QN(n5748) );
  DFFRX1 \CACHE_reg[3][66]  ( .D(n4509), .CK(clk), .RN(n3053), .Q(
        \CACHE[3][66] ), .QN(n5749) );
  DFFRX1 \CACHE_reg[3][65]  ( .D(n4510), .CK(clk), .RN(n3054), .Q(
        \CACHE[3][65] ), .QN(n5750) );
  DFFRX1 \CACHE_reg[3][64]  ( .D(n4511), .CK(clk), .RN(n3054), .Q(
        \CACHE[3][64] ), .QN(n5751) );
  DFFRX1 \CACHE_reg[3][63]  ( .D(n4512), .CK(clk), .RN(n512), .Q(
        \CACHE[3][63] ), .QN(n5752) );
  DFFRX1 \CACHE_reg[3][62]  ( .D(n4513), .CK(clk), .RN(n513), .Q(
        \CACHE[3][62] ), .QN(n5753) );
  DFFRX1 \CACHE_reg[3][61]  ( .D(n4514), .CK(clk), .RN(n514), .Q(
        \CACHE[3][61] ), .QN(n5754) );
  DFFRX1 \CACHE_reg[3][60]  ( .D(n4515), .CK(clk), .RN(n514), .Q(
        \CACHE[3][60] ), .QN(n5755) );
  DFFRX1 \CACHE_reg[3][59]  ( .D(n4516), .CK(clk), .RN(n515), .Q(
        \CACHE[3][59] ), .QN(n5756) );
  DFFRX1 \CACHE_reg[3][58]  ( .D(n4517), .CK(clk), .RN(n516), .Q(
        \CACHE[3][58] ), .QN(n5757) );
  DFFRX1 \CACHE_reg[3][57]  ( .D(n4518), .CK(clk), .RN(n516), .Q(
        \CACHE[3][57] ), .QN(n5758) );
  DFFRX1 \CACHE_reg[3][56]  ( .D(n4519), .CK(clk), .RN(n517), .Q(
        \CACHE[3][56] ), .QN(n5759) );
  DFFRX1 \CACHE_reg[3][55]  ( .D(n4520), .CK(clk), .RN(n518), .Q(
        \CACHE[3][55] ), .QN(n5760) );
  DFFRX1 \CACHE_reg[3][54]  ( .D(n4521), .CK(clk), .RN(n518), .Q(
        \CACHE[3][54] ), .QN(n5761) );
  DFFRX1 \CACHE_reg[3][53]  ( .D(n4522), .CK(clk), .RN(n519), .Q(
        \CACHE[3][53] ), .QN(n5762) );
  DFFRX1 \CACHE_reg[3][52]  ( .D(n4523), .CK(clk), .RN(n520), .Q(
        \CACHE[3][52] ), .QN(n5763) );
  DFFRX1 \CACHE_reg[3][51]  ( .D(n4524), .CK(clk), .RN(n520), .Q(
        \CACHE[3][51] ), .QN(n5764) );
  DFFRX1 \CACHE_reg[3][50]  ( .D(n4525), .CK(clk), .RN(n521), .Q(
        \CACHE[3][50] ), .QN(n5765) );
  DFFRX1 \CACHE_reg[3][49]  ( .D(n4526), .CK(clk), .RN(n522), .Q(
        \CACHE[3][49] ), .QN(n5766) );
  DFFRX1 \CACHE_reg[3][48]  ( .D(n4527), .CK(clk), .RN(n522), .Q(
        \CACHE[3][48] ), .QN(n5767) );
  DFFRX1 \CACHE_reg[3][47]  ( .D(n4528), .CK(clk), .RN(n523), .Q(
        \CACHE[3][47] ), .QN(n5768) );
  DFFRX1 \CACHE_reg[3][46]  ( .D(n4529), .CK(clk), .RN(n524), .Q(
        \CACHE[3][46] ), .QN(n5769) );
  DFFRX1 \CACHE_reg[3][45]  ( .D(n4530), .CK(clk), .RN(n524), .Q(
        \CACHE[3][45] ), .QN(n5770) );
  DFFRX1 \CACHE_reg[3][44]  ( .D(n4531), .CK(clk), .RN(n525), .Q(
        \CACHE[3][44] ), .QN(n5771) );
  DFFRX1 \CACHE_reg[3][43]  ( .D(n4532), .CK(clk), .RN(n526), .Q(
        \CACHE[3][43] ), .QN(n5772) );
  DFFRX1 \CACHE_reg[3][42]  ( .D(n4533), .CK(clk), .RN(n526), .Q(
        \CACHE[3][42] ), .QN(n5773) );
  DFFRX1 \CACHE_reg[3][41]  ( .D(n4534), .CK(clk), .RN(n527), .Q(
        \CACHE[3][41] ), .QN(n5774) );
  DFFRX1 \CACHE_reg[3][40]  ( .D(n4535), .CK(clk), .RN(n528), .Q(
        \CACHE[3][40] ), .QN(n5775) );
  DFFRX1 \CACHE_reg[3][39]  ( .D(n4536), .CK(clk), .RN(n528), .Q(
        \CACHE[3][39] ), .QN(n5776) );
  DFFRX1 \CACHE_reg[3][38]  ( .D(n4537), .CK(clk), .RN(n529), .Q(
        \CACHE[3][38] ), .QN(n5777) );
  DFFRX1 \CACHE_reg[3][37]  ( .D(n4538), .CK(clk), .RN(n530), .Q(
        \CACHE[3][37] ), .QN(n5778) );
  DFFRX1 \CACHE_reg[3][36]  ( .D(n4539), .CK(clk), .RN(n530), .Q(
        \CACHE[3][36] ), .QN(n5779) );
  DFFRX1 \CACHE_reg[3][35]  ( .D(n4540), .CK(clk), .RN(n531), .Q(
        \CACHE[3][35] ), .QN(n5780) );
  DFFRX1 \CACHE_reg[3][34]  ( .D(n4541), .CK(clk), .RN(n532), .Q(
        \CACHE[3][34] ), .QN(n5781) );
  DFFRX1 \CACHE_reg[3][33]  ( .D(n4542), .CK(clk), .RN(n532), .Q(
        \CACHE[3][33] ), .QN(n5782) );
  DFFRX1 \CACHE_reg[3][32]  ( .D(n4543), .CK(clk), .RN(n533), .Q(
        \CACHE[3][32] ), .QN(n5783) );
  DFFRX1 \CACHE_reg[3][31]  ( .D(n4544), .CK(clk), .RN(n491), .Q(
        \CACHE[3][31] ), .QN(n5784) );
  DFFRX1 \CACHE_reg[3][30]  ( .D(n4545), .CK(clk), .RN(n3055), .Q(
        \CACHE[3][30] ), .QN(n5785) );
  DFFRX1 \CACHE_reg[3][29]  ( .D(n4546), .CK(clk), .RN(n492), .Q(
        \CACHE[3][29] ), .QN(n5786) );
  DFFRX1 \CACHE_reg[3][28]  ( .D(n4547), .CK(clk), .RN(n493), .Q(
        \CACHE[3][28] ), .QN(n5787) );
  DFFRX1 \CACHE_reg[3][27]  ( .D(n4548), .CK(clk), .RN(n494), .Q(
        \CACHE[3][27] ), .QN(n5788) );
  DFFRX1 \CACHE_reg[3][26]  ( .D(n4549), .CK(clk), .RN(n494), .Q(
        \CACHE[3][26] ), .QN(n5789) );
  DFFRX1 \CACHE_reg[3][25]  ( .D(n4550), .CK(clk), .RN(n495), .Q(
        \CACHE[3][25] ), .QN(n5790) );
  DFFRX1 \CACHE_reg[3][24]  ( .D(n4551), .CK(clk), .RN(n496), .Q(
        \CACHE[3][24] ), .QN(n5791) );
  DFFRX1 \CACHE_reg[3][23]  ( .D(n4552), .CK(clk), .RN(n496), .Q(
        \CACHE[3][23] ), .QN(n5792) );
  DFFRX1 \CACHE_reg[3][22]  ( .D(n4553), .CK(clk), .RN(n497), .Q(
        \CACHE[3][22] ), .QN(n5793) );
  DFFRX1 \CACHE_reg[3][21]  ( .D(n4554), .CK(clk), .RN(n498), .Q(
        \CACHE[3][21] ), .QN(n5794) );
  DFFRX1 \CACHE_reg[3][20]  ( .D(n4555), .CK(clk), .RN(n498), .Q(
        \CACHE[3][20] ), .QN(n5795) );
  DFFRX1 \CACHE_reg[3][19]  ( .D(n4556), .CK(clk), .RN(n499), .Q(
        \CACHE[3][19] ), .QN(n5796) );
  DFFRX1 \CACHE_reg[3][18]  ( .D(n4557), .CK(clk), .RN(n500), .Q(
        \CACHE[3][18] ), .QN(n5797) );
  DFFRX1 \CACHE_reg[3][17]  ( .D(n4558), .CK(clk), .RN(n500), .Q(
        \CACHE[3][17] ), .QN(n5798) );
  DFFRX1 \CACHE_reg[3][16]  ( .D(n4559), .CK(clk), .RN(n501), .Q(
        \CACHE[3][16] ), .QN(n5799) );
  DFFRX1 \CACHE_reg[3][15]  ( .D(n4560), .CK(clk), .RN(n502), .Q(
        \CACHE[3][15] ), .QN(n5800) );
  DFFRX1 \CACHE_reg[3][14]  ( .D(n4561), .CK(clk), .RN(n502), .Q(
        \CACHE[3][14] ), .QN(n5801) );
  DFFRX1 \CACHE_reg[3][13]  ( .D(n4562), .CK(clk), .RN(n503), .Q(
        \CACHE[3][13] ), .QN(n5802) );
  DFFRX1 \CACHE_reg[3][12]  ( .D(n4563), .CK(clk), .RN(n504), .Q(
        \CACHE[3][12] ), .QN(n5803) );
  DFFRX1 \CACHE_reg[3][11]  ( .D(n4564), .CK(clk), .RN(n504), .Q(
        \CACHE[3][11] ), .QN(n5804) );
  DFFRX1 \CACHE_reg[3][10]  ( .D(n4565), .CK(clk), .RN(n505), .Q(
        \CACHE[3][10] ), .QN(n5805) );
  DFFRX1 \CACHE_reg[3][9]  ( .D(n4566), .CK(clk), .RN(n506), .Q(\CACHE[3][9] ), 
        .QN(n5806) );
  DFFRX1 \CACHE_reg[3][8]  ( .D(n4567), .CK(clk), .RN(n506), .Q(\CACHE[3][8] ), 
        .QN(n5807) );
  DFFRX1 \CACHE_reg[3][7]  ( .D(n4568), .CK(clk), .RN(n507), .Q(\CACHE[3][7] ), 
        .QN(n5808) );
  DFFRX1 \CACHE_reg[3][6]  ( .D(n4569), .CK(clk), .RN(n508), .Q(\CACHE[3][6] ), 
        .QN(n5809) );
  DFFRX1 \CACHE_reg[3][5]  ( .D(n4570), .CK(clk), .RN(n508), .Q(\CACHE[3][5] ), 
        .QN(n5810) );
  DFFRX1 \CACHE_reg[3][4]  ( .D(n4571), .CK(clk), .RN(n509), .Q(\CACHE[3][4] ), 
        .QN(n5811) );
  DFFRX1 \CACHE_reg[3][3]  ( .D(n4572), .CK(clk), .RN(n510), .Q(\CACHE[3][3] ), 
        .QN(n5812) );
  DFFRX1 \CACHE_reg[3][2]  ( .D(n4573), .CK(clk), .RN(n510), .Q(\CACHE[3][2] ), 
        .QN(n5813) );
  DFFRX1 \CACHE_reg[3][1]  ( .D(n4574), .CK(clk), .RN(n511), .Q(\CACHE[3][1] ), 
        .QN(n5814) );
  DFFRX1 \CACHE_reg[3][0]  ( .D(n4575), .CK(clk), .RN(n512), .Q(\CACHE[3][0] ), 
        .QN(n5815) );
  DFFRX1 \CACHE_reg[5][154]  ( .D(n4111), .CK(clk), .RN(n492), .Q(
        \CACHE[5][154] ), .QN(n5351) );
  DFFRX1 \CACHE_reg[5][153]  ( .D(n4112), .CK(clk), .RN(n492), .Q(
        \CACHE[5][153] ), .QN(n5352) );
  DFFRX1 \CACHE_reg[5][152]  ( .D(n4113), .CK(clk), .RN(n474), .Q(
        \CACHE[5][152] ), .QN(n5353) );
  DFFRX1 \CACHE_reg[5][151]  ( .D(n4114), .CK(clk), .RN(n475), .Q(
        \CACHE[5][151] ), .QN(n5354) );
  DFFRX1 \CACHE_reg[5][150]  ( .D(n4115), .CK(clk), .RN(n476), .Q(
        \CACHE[5][150] ), .QN(n5355) );
  DFFRX1 \CACHE_reg[5][149]  ( .D(n4116), .CK(clk), .RN(n476), .Q(
        \CACHE[5][149] ), .QN(n5356) );
  DFFRX1 \CACHE_reg[5][148]  ( .D(n4117), .CK(clk), .RN(n477), .Q(
        \CACHE[5][148] ), .QN(n5357) );
  DFFRX1 \CACHE_reg[5][147]  ( .D(n4118), .CK(clk), .RN(n478), .Q(
        \CACHE[5][147] ), .QN(n5358) );
  DFFRX1 \CACHE_reg[5][146]  ( .D(n4119), .CK(clk), .RN(n478), .Q(
        \CACHE[5][146] ), .QN(n5359) );
  DFFRX1 \CACHE_reg[5][145]  ( .D(n4120), .CK(clk), .RN(n479), .Q(
        \CACHE[5][145] ), .QN(n5360) );
  DFFRX1 \CACHE_reg[5][144]  ( .D(n4121), .CK(clk), .RN(n480), .Q(
        \CACHE[5][144] ), .QN(n5361) );
  DFFRX1 \CACHE_reg[5][143]  ( .D(n4122), .CK(clk), .RN(n480), .Q(
        \CACHE[5][143] ), .QN(n5362) );
  DFFRX1 \CACHE_reg[5][142]  ( .D(n4123), .CK(clk), .RN(n481), .Q(
        \CACHE[5][142] ), .QN(n5363) );
  DFFRX1 \CACHE_reg[5][141]  ( .D(n4124), .CK(clk), .RN(n482), .Q(
        \CACHE[5][141] ), .QN(n5364) );
  DFFRX1 \CACHE_reg[5][140]  ( .D(n4125), .CK(clk), .RN(n482), .Q(
        \CACHE[5][140] ), .QN(n5365) );
  DFFRX1 \CACHE_reg[5][139]  ( .D(n4126), .CK(clk), .RN(n490), .Q(
        \CACHE[5][139] ), .QN(n5366) );
  DFFRX1 \CACHE_reg[5][138]  ( .D(n4127), .CK(clk), .RN(n483), .Q(
        \CACHE[5][138] ), .QN(n5367) );
  DFFRX1 \CACHE_reg[5][137]  ( .D(n4128), .CK(clk), .RN(n484), .Q(
        \CACHE[5][137] ), .QN(n5368) );
  DFFRX1 \CACHE_reg[5][136]  ( .D(n4129), .CK(clk), .RN(n484), .Q(
        \CACHE[5][136] ), .QN(n5369) );
  DFFRX1 \CACHE_reg[5][135]  ( .D(n4130), .CK(clk), .RN(n485), .Q(
        \CACHE[5][135] ), .QN(n5370) );
  DFFRX1 \CACHE_reg[5][134]  ( .D(n4131), .CK(clk), .RN(n486), .Q(
        \CACHE[5][134] ), .QN(n5371) );
  DFFRX1 \CACHE_reg[5][133]  ( .D(n4132), .CK(clk), .RN(n486), .Q(
        \CACHE[5][133] ), .QN(n5372) );
  DFFRX1 \CACHE_reg[5][132]  ( .D(n4133), .CK(clk), .RN(n474), .Q(
        \CACHE[5][132] ), .QN(n5373) );
  DFFRX1 \CACHE_reg[5][131]  ( .D(n4134), .CK(clk), .RN(n487), .Q(
        \CACHE[5][131] ), .QN(n5374) );
  DFFRX1 \CACHE_reg[5][130]  ( .D(n4135), .CK(clk), .RN(n488), .Q(
        \CACHE[5][130] ), .QN(n5375) );
  DFFRX1 \CACHE_reg[5][129]  ( .D(n4136), .CK(clk), .RN(n488), .Q(
        \CACHE[5][129] ), .QN(n5376) );
  DFFRX1 \CACHE_reg[5][128]  ( .D(n4137), .CK(clk), .RN(n489), .Q(
        \CACHE[5][128] ), .QN(n5377) );
  DFFRX1 \CACHE_reg[5][127]  ( .D(n4138), .CK(clk), .RN(n492), .Q(
        \CACHE[5][127] ), .QN(n5378) );
  DFFRX1 \CACHE_reg[5][126]  ( .D(n4139), .CK(clk), .RN(n491), .Q(
        \CACHE[5][126] ), .QN(n5379) );
  DFFRX1 \CACHE_reg[5][125]  ( .D(n4140), .CK(clk), .RN(n492), .Q(
        \CACHE[5][125] ), .QN(n5380) );
  DFFRX1 \CACHE_reg[5][124]  ( .D(n4141), .CK(clk), .RN(n3055), .Q(
        \CACHE[5][124] ), .QN(n5381) );
  DFFRX1 \CACHE_reg[5][123]  ( .D(n4142), .CK(clk), .RN(n535), .Q(
        \CACHE[5][123] ), .QN(n5382) );
  DFFRX1 \CACHE_reg[5][122]  ( .D(n4143), .CK(clk), .RN(n535), .Q(
        \CACHE[5][122] ), .QN(n5383) );
  DFFRX1 \CACHE_reg[5][121]  ( .D(n4144), .CK(clk), .RN(n536), .Q(
        \CACHE[5][121] ), .QN(n5384) );
  DFFRX1 \CACHE_reg[5][120]  ( .D(n4145), .CK(clk), .RN(n537), .Q(
        \CACHE[5][120] ), .QN(n5385) );
  DFFRX1 \CACHE_reg[5][119]  ( .D(n4146), .CK(clk), .RN(n537), .Q(
        \CACHE[5][119] ), .QN(n5386) );
  DFFRX1 \CACHE_reg[5][118]  ( .D(n4147), .CK(clk), .RN(n538), .Q(
        \CACHE[5][118] ), .QN(n5387) );
  DFFRX1 \CACHE_reg[5][117]  ( .D(n4148), .CK(clk), .RN(n539), .Q(
        \CACHE[5][117] ), .QN(n5388) );
  DFFRX1 \CACHE_reg[5][116]  ( .D(n4149), .CK(clk), .RN(n539), .Q(
        \CACHE[5][116] ), .QN(n5389) );
  DFFRX1 \CACHE_reg[5][115]  ( .D(n4150), .CK(clk), .RN(n540), .Q(
        \CACHE[5][115] ), .QN(n5390) );
  DFFRX1 \CACHE_reg[5][114]  ( .D(n4151), .CK(clk), .RN(n3020), .Q(
        \CACHE[5][114] ), .QN(n5391) );
  DFFRX1 \CACHE_reg[5][113]  ( .D(n4152), .CK(clk), .RN(n3020), .Q(
        \CACHE[5][113] ), .QN(n5392) );
  DFFRX1 \CACHE_reg[5][112]  ( .D(n4153), .CK(clk), .RN(n3022), .Q(
        \CACHE[5][112] ), .QN(n5393) );
  DFFRX1 \CACHE_reg[5][111]  ( .D(n4154), .CK(clk), .RN(n3023), .Q(
        \CACHE[5][111] ), .QN(n5394) );
  DFFRX1 \CACHE_reg[5][110]  ( .D(n4155), .CK(clk), .RN(n3023), .Q(
        \CACHE[5][110] ), .QN(n5395) );
  DFFRX1 \CACHE_reg[5][109]  ( .D(n4156), .CK(clk), .RN(n3024), .Q(
        \CACHE[5][109] ), .QN(n5396) );
  DFFRX1 \CACHE_reg[5][108]  ( .D(n4157), .CK(clk), .RN(n3025), .Q(
        \CACHE[5][108] ), .QN(n5397) );
  DFFRX1 \CACHE_reg[5][107]  ( .D(n4158), .CK(clk), .RN(n3025), .Q(
        \CACHE[5][107] ), .QN(n5398) );
  DFFRX1 \CACHE_reg[5][106]  ( .D(n4159), .CK(clk), .RN(n3026), .Q(
        \CACHE[5][106] ), .QN(n5399) );
  DFFRX1 \CACHE_reg[5][105]  ( .D(n4160), .CK(clk), .RN(n3027), .Q(
        \CACHE[5][105] ), .QN(n5400) );
  DFFRX1 \CACHE_reg[5][104]  ( .D(n4161), .CK(clk), .RN(n3027), .Q(
        \CACHE[5][104] ), .QN(n5401) );
  DFFRX1 \CACHE_reg[5][103]  ( .D(n4162), .CK(clk), .RN(n3028), .Q(
        \CACHE[5][103] ), .QN(n5402) );
  DFFRX1 \CACHE_reg[5][102]  ( .D(n4163), .CK(clk), .RN(n3029), .Q(
        \CACHE[5][102] ), .QN(n5403) );
  DFFRX1 \CACHE_reg[5][101]  ( .D(n4164), .CK(clk), .RN(n3029), .Q(
        \CACHE[5][101] ), .QN(n5404) );
  DFFRX1 \CACHE_reg[5][100]  ( .D(n4165), .CK(clk), .RN(n3030), .Q(
        \CACHE[5][100] ), .QN(n5405) );
  DFFRX1 \CACHE_reg[5][99]  ( .D(n4166), .CK(clk), .RN(n3031), .Q(
        \CACHE[5][99] ), .QN(n5406) );
  DFFRX1 \CACHE_reg[5][98]  ( .D(n4167), .CK(clk), .RN(n3031), .Q(
        \CACHE[5][98] ), .QN(n5407) );
  DFFRX1 \CACHE_reg[5][97]  ( .D(n4168), .CK(clk), .RN(n3032), .Q(
        \CACHE[5][97] ), .QN(n5408) );
  DFFRX1 \CACHE_reg[5][96]  ( .D(n4169), .CK(clk), .RN(n3033), .Q(
        \CACHE[5][96] ), .QN(n5409) );
  DFFRX1 \CACHE_reg[5][95]  ( .D(n4170), .CK(clk), .RN(n3033), .Q(
        \CACHE[5][95] ), .QN(n5410) );
  DFFRX1 \CACHE_reg[5][94]  ( .D(n4171), .CK(clk), .RN(n3034), .Q(
        \CACHE[5][94] ), .QN(n5411) );
  DFFRX1 \CACHE_reg[5][93]  ( .D(n4172), .CK(clk), .RN(n3035), .Q(
        \CACHE[5][93] ), .QN(n5412) );
  DFFRX1 \CACHE_reg[5][92]  ( .D(n4173), .CK(clk), .RN(n3035), .Q(
        \CACHE[5][92] ), .QN(n5413) );
  DFFRX1 \CACHE_reg[5][91]  ( .D(n4174), .CK(clk), .RN(n3036), .Q(
        \CACHE[5][91] ), .QN(n5414) );
  DFFRX1 \CACHE_reg[5][90]  ( .D(n4175), .CK(clk), .RN(n3037), .Q(
        \CACHE[5][90] ), .QN(n5415) );
  DFFRX1 \CACHE_reg[5][89]  ( .D(n4176), .CK(clk), .RN(n3037), .Q(
        \CACHE[5][89] ), .QN(n5416) );
  DFFRX1 \CACHE_reg[5][88]  ( .D(n4177), .CK(clk), .RN(n3038), .Q(
        \CACHE[5][88] ), .QN(n5417) );
  DFFRX1 \CACHE_reg[5][87]  ( .D(n4178), .CK(clk), .RN(n3039), .Q(
        \CACHE[5][87] ), .QN(n5418) );
  DFFRX1 \CACHE_reg[5][86]  ( .D(n4179), .CK(clk), .RN(n3039), .Q(
        \CACHE[5][86] ), .QN(n5419) );
  DFFRX1 \CACHE_reg[5][85]  ( .D(n4180), .CK(clk), .RN(n3040), .Q(
        \CACHE[5][85] ), .QN(n5420) );
  DFFRX1 \CACHE_reg[5][84]  ( .D(n4181), .CK(clk), .RN(n3041), .Q(
        \CACHE[5][84] ), .QN(n5421) );
  DFFRX1 \CACHE_reg[5][83]  ( .D(n4182), .CK(clk), .RN(n3041), .Q(
        \CACHE[5][83] ), .QN(n5422) );
  DFFRX1 \CACHE_reg[5][82]  ( .D(n4183), .CK(clk), .RN(n3042), .Q(
        \CACHE[5][82] ), .QN(n5423) );
  DFFRX1 \CACHE_reg[5][81]  ( .D(n4184), .CK(clk), .RN(n3043), .Q(
        \CACHE[5][81] ), .QN(n5424) );
  DFFRX1 \CACHE_reg[5][80]  ( .D(n4185), .CK(clk), .RN(n3043), .Q(
        \CACHE[5][80] ), .QN(n5425) );
  DFFRX1 \CACHE_reg[5][79]  ( .D(n4186), .CK(clk), .RN(n3044), .Q(
        \CACHE[5][79] ), .QN(n5426) );
  DFFRX1 \CACHE_reg[5][78]  ( .D(n4187), .CK(clk), .RN(n3045), .Q(
        \CACHE[5][78] ), .QN(n5427) );
  DFFRX1 \CACHE_reg[5][77]  ( .D(n4188), .CK(clk), .RN(n3045), .Q(
        \CACHE[5][77] ), .QN(n5428) );
  DFFRX1 \CACHE_reg[5][76]  ( .D(n4189), .CK(clk), .RN(n3046), .Q(
        \CACHE[5][76] ), .QN(n5429) );
  DFFRX1 \CACHE_reg[5][75]  ( .D(n4190), .CK(clk), .RN(n3047), .Q(
        \CACHE[5][75] ), .QN(n5430) );
  DFFRX1 \CACHE_reg[5][74]  ( .D(n4191), .CK(clk), .RN(n3047), .Q(
        \CACHE[5][74] ), .QN(n5431) );
  DFFRX1 \CACHE_reg[5][73]  ( .D(n4192), .CK(clk), .RN(n3048), .Q(
        \CACHE[5][73] ), .QN(n5432) );
  DFFRX1 \CACHE_reg[5][72]  ( .D(n4193), .CK(clk), .RN(n3049), .Q(
        \CACHE[5][72] ), .QN(n5433) );
  DFFRX1 \CACHE_reg[5][71]  ( .D(n4194), .CK(clk), .RN(n3049), .Q(
        \CACHE[5][71] ), .QN(n5434) );
  DFFRX1 \CACHE_reg[5][70]  ( .D(n4195), .CK(clk), .RN(n3050), .Q(
        \CACHE[5][70] ), .QN(n5435) );
  DFFRX1 \CACHE_reg[5][69]  ( .D(n4196), .CK(clk), .RN(n3051), .Q(
        \CACHE[5][69] ), .QN(n5436) );
  DFFRX1 \CACHE_reg[5][68]  ( .D(n4197), .CK(clk), .RN(n3051), .Q(
        \CACHE[5][68] ), .QN(n5437) );
  DFFRX1 \CACHE_reg[5][67]  ( .D(n4198), .CK(clk), .RN(n3052), .Q(
        \CACHE[5][67] ), .QN(n5438) );
  DFFRX1 \CACHE_reg[5][66]  ( .D(n4199), .CK(clk), .RN(n3053), .Q(
        \CACHE[5][66] ), .QN(n5439) );
  DFFRX1 \CACHE_reg[5][65]  ( .D(n4200), .CK(clk), .RN(n3053), .Q(
        \CACHE[5][65] ), .QN(n5440) );
  DFFRX1 \CACHE_reg[5][64]  ( .D(n4201), .CK(clk), .RN(n3054), .Q(
        \CACHE[5][64] ), .QN(n5441) );
  DFFRX1 \CACHE_reg[5][63]  ( .D(n4202), .CK(clk), .RN(n512), .Q(
        \CACHE[5][63] ), .QN(n5442) );
  DFFRX1 \CACHE_reg[5][62]  ( .D(n4203), .CK(clk), .RN(n513), .Q(
        \CACHE[5][62] ), .QN(n5443) );
  DFFRX1 \CACHE_reg[5][61]  ( .D(n4204), .CK(clk), .RN(n514), .Q(
        \CACHE[5][61] ), .QN(n5444) );
  DFFRX1 \CACHE_reg[5][60]  ( .D(n4205), .CK(clk), .RN(n514), .Q(
        \CACHE[5][60] ), .QN(n5445) );
  DFFRX1 \CACHE_reg[5][59]  ( .D(n4206), .CK(clk), .RN(n515), .Q(
        \CACHE[5][59] ), .QN(n5446) );
  DFFRX1 \CACHE_reg[5][58]  ( .D(n4207), .CK(clk), .RN(n516), .Q(
        \CACHE[5][58] ), .QN(n5447) );
  DFFRX1 \CACHE_reg[5][57]  ( .D(n4208), .CK(clk), .RN(n516), .Q(
        \CACHE[5][57] ), .QN(n5448) );
  DFFRX1 \CACHE_reg[5][56]  ( .D(n4209), .CK(clk), .RN(n517), .Q(
        \CACHE[5][56] ), .QN(n5449) );
  DFFRX1 \CACHE_reg[5][55]  ( .D(n4210), .CK(clk), .RN(n518), .Q(
        \CACHE[5][55] ), .QN(n5450) );
  DFFRX1 \CACHE_reg[5][54]  ( .D(n4211), .CK(clk), .RN(n518), .Q(
        \CACHE[5][54] ), .QN(n5451) );
  DFFRX1 \CACHE_reg[5][53]  ( .D(n4212), .CK(clk), .RN(n519), .Q(
        \CACHE[5][53] ), .QN(n5452) );
  DFFRX1 \CACHE_reg[5][52]  ( .D(n4213), .CK(clk), .RN(n520), .Q(
        \CACHE[5][52] ), .QN(n5453) );
  DFFRX1 \CACHE_reg[5][51]  ( .D(n4214), .CK(clk), .RN(n520), .Q(
        \CACHE[5][51] ), .QN(n5454) );
  DFFRX1 \CACHE_reg[5][50]  ( .D(n4215), .CK(clk), .RN(n521), .Q(
        \CACHE[5][50] ), .QN(n5455) );
  DFFRX1 \CACHE_reg[5][49]  ( .D(n4216), .CK(clk), .RN(n522), .Q(
        \CACHE[5][49] ), .QN(n5456) );
  DFFRX1 \CACHE_reg[5][48]  ( .D(n4217), .CK(clk), .RN(n522), .Q(
        \CACHE[5][48] ), .QN(n5457) );
  DFFRX1 \CACHE_reg[5][47]  ( .D(n4218), .CK(clk), .RN(n523), .Q(
        \CACHE[5][47] ), .QN(n5458) );
  DFFRX1 \CACHE_reg[5][46]  ( .D(n4219), .CK(clk), .RN(n524), .Q(
        \CACHE[5][46] ), .QN(n5459) );
  DFFRX1 \CACHE_reg[5][45]  ( .D(n4220), .CK(clk), .RN(n524), .Q(
        \CACHE[5][45] ), .QN(n5460) );
  DFFRX1 \CACHE_reg[5][44]  ( .D(n4221), .CK(clk), .RN(n525), .Q(
        \CACHE[5][44] ), .QN(n5461) );
  DFFRX1 \CACHE_reg[5][43]  ( .D(n4222), .CK(clk), .RN(n526), .Q(
        \CACHE[5][43] ), .QN(n5462) );
  DFFRX1 \CACHE_reg[5][42]  ( .D(n4223), .CK(clk), .RN(n526), .Q(
        \CACHE[5][42] ), .QN(n5463) );
  DFFRX1 \CACHE_reg[5][41]  ( .D(n4224), .CK(clk), .RN(n527), .Q(
        \CACHE[5][41] ), .QN(n5464) );
  DFFRX1 \CACHE_reg[5][40]  ( .D(n4225), .CK(clk), .RN(n528), .Q(
        \CACHE[5][40] ), .QN(n5465) );
  DFFRX1 \CACHE_reg[5][39]  ( .D(n4226), .CK(clk), .RN(n528), .Q(
        \CACHE[5][39] ), .QN(n5466) );
  DFFRX1 \CACHE_reg[5][38]  ( .D(n4227), .CK(clk), .RN(n529), .Q(
        \CACHE[5][38] ), .QN(n5467) );
  DFFRX1 \CACHE_reg[5][37]  ( .D(n4228), .CK(clk), .RN(n530), .Q(
        \CACHE[5][37] ), .QN(n5468) );
  DFFRX1 \CACHE_reg[5][36]  ( .D(n4229), .CK(clk), .RN(n530), .Q(
        \CACHE[5][36] ), .QN(n5469) );
  DFFRX1 \CACHE_reg[5][35]  ( .D(n4230), .CK(clk), .RN(n531), .Q(
        \CACHE[5][35] ), .QN(n5470) );
  DFFRX1 \CACHE_reg[5][34]  ( .D(n4231), .CK(clk), .RN(n532), .Q(
        \CACHE[5][34] ), .QN(n5471) );
  DFFRX1 \CACHE_reg[5][33]  ( .D(n4232), .CK(clk), .RN(n532), .Q(
        \CACHE[5][33] ), .QN(n5472) );
  DFFRX1 \CACHE_reg[5][32]  ( .D(n4233), .CK(clk), .RN(n533), .Q(
        \CACHE[5][32] ), .QN(n5473) );
  DFFRX1 \CACHE_reg[5][31]  ( .D(n4234), .CK(clk), .RN(n490), .Q(
        \CACHE[5][31] ), .QN(n5474) );
  DFFRX1 \CACHE_reg[5][30]  ( .D(n4235), .CK(clk), .RN(n3055), .Q(
        \CACHE[5][30] ), .QN(n5475) );
  DFFRX1 \CACHE_reg[5][29]  ( .D(n4236), .CK(clk), .RN(n492), .Q(
        \CACHE[5][29] ), .QN(n5476) );
  DFFRX1 \CACHE_reg[5][28]  ( .D(n4237), .CK(clk), .RN(n493), .Q(
        \CACHE[5][28] ), .QN(n5477) );
  DFFRX1 \CACHE_reg[5][27]  ( .D(n4238), .CK(clk), .RN(n494), .Q(
        \CACHE[5][27] ), .QN(n5478) );
  DFFRX1 \CACHE_reg[5][26]  ( .D(n4239), .CK(clk), .RN(n494), .Q(
        \CACHE[5][26] ), .QN(n5479) );
  DFFRX1 \CACHE_reg[5][25]  ( .D(n4240), .CK(clk), .RN(n495), .Q(
        \CACHE[5][25] ), .QN(n5480) );
  DFFRX1 \CACHE_reg[5][24]  ( .D(n4241), .CK(clk), .RN(n496), .Q(
        \CACHE[5][24] ), .QN(n5481) );
  DFFRX1 \CACHE_reg[5][23]  ( .D(n4242), .CK(clk), .RN(n496), .Q(
        \CACHE[5][23] ), .QN(n5482) );
  DFFRX1 \CACHE_reg[5][22]  ( .D(n4243), .CK(clk), .RN(n497), .Q(
        \CACHE[5][22] ), .QN(n5483) );
  DFFRX1 \CACHE_reg[5][21]  ( .D(n4244), .CK(clk), .RN(n498), .Q(
        \CACHE[5][21] ), .QN(n5484) );
  DFFRX1 \CACHE_reg[5][20]  ( .D(n4245), .CK(clk), .RN(n498), .Q(
        \CACHE[5][20] ), .QN(n5485) );
  DFFRX1 \CACHE_reg[5][19]  ( .D(n4246), .CK(clk), .RN(n499), .Q(
        \CACHE[5][19] ), .QN(n5486) );
  DFFRX1 \CACHE_reg[5][18]  ( .D(n4247), .CK(clk), .RN(n500), .Q(
        \CACHE[5][18] ), .QN(n5487) );
  DFFRX1 \CACHE_reg[5][17]  ( .D(n4248), .CK(clk), .RN(n500), .Q(
        \CACHE[5][17] ), .QN(n5488) );
  DFFRX1 \CACHE_reg[5][16]  ( .D(n4249), .CK(clk), .RN(n501), .Q(
        \CACHE[5][16] ), .QN(n5489) );
  DFFRX1 \CACHE_reg[5][15]  ( .D(n4250), .CK(clk), .RN(n502), .Q(
        \CACHE[5][15] ), .QN(n5490) );
  DFFRX1 \CACHE_reg[5][14]  ( .D(n4251), .CK(clk), .RN(n502), .Q(
        \CACHE[5][14] ), .QN(n5491) );
  DFFRX1 \CACHE_reg[5][13]  ( .D(n4252), .CK(clk), .RN(n503), .Q(
        \CACHE[5][13] ), .QN(n5492) );
  DFFRX1 \CACHE_reg[5][12]  ( .D(n4253), .CK(clk), .RN(n504), .Q(
        \CACHE[5][12] ), .QN(n5493) );
  DFFRX1 \CACHE_reg[5][11]  ( .D(n4254), .CK(clk), .RN(n504), .Q(
        \CACHE[5][11] ), .QN(n5494) );
  DFFRX1 \CACHE_reg[5][10]  ( .D(n4255), .CK(clk), .RN(n505), .Q(
        \CACHE[5][10] ), .QN(n5495) );
  DFFRX1 \CACHE_reg[5][9]  ( .D(n4256), .CK(clk), .RN(n506), .Q(\CACHE[5][9] ), 
        .QN(n5496) );
  DFFRX1 \CACHE_reg[5][8]  ( .D(n4257), .CK(clk), .RN(n506), .Q(\CACHE[5][8] ), 
        .QN(n5497) );
  DFFRX1 \CACHE_reg[5][7]  ( .D(n4258), .CK(clk), .RN(n507), .Q(\CACHE[5][7] ), 
        .QN(n5498) );
  DFFRX1 \CACHE_reg[5][6]  ( .D(n4259), .CK(clk), .RN(n508), .Q(\CACHE[5][6] ), 
        .QN(n5499) );
  DFFRX1 \CACHE_reg[5][5]  ( .D(n4260), .CK(clk), .RN(n508), .Q(\CACHE[5][5] ), 
        .QN(n5500) );
  DFFRX1 \CACHE_reg[5][4]  ( .D(n4261), .CK(clk), .RN(n509), .Q(\CACHE[5][4] ), 
        .QN(n5501) );
  DFFRX1 \CACHE_reg[5][3]  ( .D(n4262), .CK(clk), .RN(n510), .Q(\CACHE[5][3] ), 
        .QN(n5502) );
  DFFRX1 \CACHE_reg[5][2]  ( .D(n4263), .CK(clk), .RN(n510), .Q(\CACHE[5][2] ), 
        .QN(n5503) );
  DFFRX1 \CACHE_reg[5][1]  ( .D(n4264), .CK(clk), .RN(n511), .Q(\CACHE[5][1] ), 
        .QN(n5504) );
  DFFRX1 \CACHE_reg[5][0]  ( .D(n4265), .CK(clk), .RN(n512), .Q(\CACHE[5][0] ), 
        .QN(n5505) );
  DFFRX1 \CACHE_reg[1][154]  ( .D(n4731), .CK(clk), .RN(n3055), .Q(
        \CACHE[1][154] ), .QN(n5971) );
  DFFRX1 \CACHE_reg[1][153]  ( .D(n4732), .CK(clk), .RN(n3055), .Q(
        \CACHE[1][153] ), .QN(n5972) );
  DFFRX1 \CACHE_reg[1][152]  ( .D(n4733), .CK(clk), .RN(n475), .Q(
        \CACHE[1][152] ), .QN(n5973) );
  DFFRX1 \CACHE_reg[1][151]  ( .D(n4734), .CK(clk), .RN(n475), .Q(
        \CACHE[1][151] ), .QN(n5974) );
  DFFRX1 \CACHE_reg[1][150]  ( .D(n4735), .CK(clk), .RN(n476), .Q(
        \CACHE[1][150] ), .QN(n5975) );
  DFFRX1 \CACHE_reg[1][149]  ( .D(n4736), .CK(clk), .RN(n477), .Q(
        \CACHE[1][149] ), .QN(n5976) );
  DFFRX1 \CACHE_reg[1][148]  ( .D(n4737), .CK(clk), .RN(n477), .Q(
        \CACHE[1][148] ), .QN(n5977) );
  DFFRX1 \CACHE_reg[1][147]  ( .D(n4738), .CK(clk), .RN(n478), .Q(
        \CACHE[1][147] ), .QN(n5978) );
  DFFRX1 \CACHE_reg[1][146]  ( .D(n4739), .CK(clk), .RN(n479), .Q(
        \CACHE[1][146] ), .QN(n5979) );
  DFFRX1 \CACHE_reg[1][145]  ( .D(n4740), .CK(clk), .RN(n479), .Q(
        \CACHE[1][145] ), .QN(n5980) );
  DFFRX1 \CACHE_reg[1][144]  ( .D(n4741), .CK(clk), .RN(n480), .Q(
        \CACHE[1][144] ), .QN(n5981) );
  DFFRX1 \CACHE_reg[1][143]  ( .D(n4742), .CK(clk), .RN(n481), .Q(
        \CACHE[1][143] ), .QN(n5982) );
  DFFRX1 \CACHE_reg[1][142]  ( .D(n4743), .CK(clk), .RN(n481), .Q(
        \CACHE[1][142] ), .QN(n5983) );
  DFFRX1 \CACHE_reg[1][141]  ( .D(n4744), .CK(clk), .RN(n482), .Q(
        \CACHE[1][141] ), .QN(n5984) );
  DFFRX1 \CACHE_reg[1][140]  ( .D(n4745), .CK(clk), .RN(n483), .Q(
        \CACHE[1][140] ), .QN(n5985) );
  DFFRX1 \CACHE_reg[1][139]  ( .D(n4746), .CK(clk), .RN(n490), .Q(
        \CACHE[1][139] ), .QN(n5986) );
  DFFRX1 \CACHE_reg[1][138]  ( .D(n4747), .CK(clk), .RN(n483), .Q(
        \CACHE[1][138] ), .QN(n5987) );
  DFFRX1 \CACHE_reg[1][137]  ( .D(n4748), .CK(clk), .RN(n484), .Q(
        \CACHE[1][137] ), .QN(n5988) );
  DFFRX1 \CACHE_reg[1][136]  ( .D(n4749), .CK(clk), .RN(n485), .Q(
        \CACHE[1][136] ), .QN(n5989) );
  DFFRX1 \CACHE_reg[1][135]  ( .D(n4750), .CK(clk), .RN(n485), .Q(
        \CACHE[1][135] ), .QN(n5990) );
  DFFRX1 \CACHE_reg[1][134]  ( .D(n4751), .CK(clk), .RN(n486), .Q(
        \CACHE[1][134] ), .QN(n5991) );
  DFFRX1 \CACHE_reg[1][133]  ( .D(n4752), .CK(clk), .RN(n487), .Q(
        \CACHE[1][133] ), .QN(n5992) );
  DFFRX1 \CACHE_reg[1][132]  ( .D(n4753), .CK(clk), .RN(n474), .Q(
        \CACHE[1][132] ), .QN(n5993) );
  DFFRX1 \CACHE_reg[1][131]  ( .D(n4754), .CK(clk), .RN(n487), .Q(
        \CACHE[1][131] ), .QN(n5994) );
  DFFRX1 \CACHE_reg[1][130]  ( .D(n4755), .CK(clk), .RN(n488), .Q(
        \CACHE[1][130] ), .QN(n5995) );
  DFFRX1 \CACHE_reg[1][129]  ( .D(n4756), .CK(clk), .RN(n489), .Q(
        \CACHE[1][129] ), .QN(n5996) );
  DFFRX1 \CACHE_reg[1][128]  ( .D(n4757), .CK(clk), .RN(n489), .Q(
        \CACHE[1][128] ), .QN(n5997) );
  DFFRX1 \CACHE_reg[1][127]  ( .D(n4758), .CK(clk), .RN(n3055), .Q(
        \CACHE[1][127] ), .QN(n5998) );
  DFFRX1 \CACHE_reg[1][126]  ( .D(n4759), .CK(clk), .RN(n492), .Q(
        \CACHE[1][126] ), .QN(n5999) );
  DFFRX1 \CACHE_reg[1][125]  ( .D(n4760), .CK(clk), .RN(n534), .Q(
        \CACHE[1][125] ), .QN(n6000) );
  DFFRX1 \CACHE_reg[1][124]  ( .D(n4761), .CK(clk), .RN(n534), .Q(
        \CACHE[1][124] ), .QN(n6001) );
  DFFRX1 \CACHE_reg[1][123]  ( .D(n4762), .CK(clk), .RN(n535), .Q(
        \CACHE[1][123] ), .QN(n6002) );
  DFFRX1 \CACHE_reg[1][122]  ( .D(n4763), .CK(clk), .RN(n536), .Q(
        \CACHE[1][122] ), .QN(n6003) );
  DFFRX1 \CACHE_reg[1][121]  ( .D(n4764), .CK(clk), .RN(n536), .Q(
        \CACHE[1][121] ), .QN(n6004) );
  DFFRX1 \CACHE_reg[1][120]  ( .D(n4765), .CK(clk), .RN(n537), .Q(
        \CACHE[1][120] ), .QN(n6005) );
  DFFRX1 \CACHE_reg[1][119]  ( .D(n4766), .CK(clk), .RN(n538), .Q(
        \CACHE[1][119] ), .QN(n6006) );
  DFFRX1 \CACHE_reg[1][118]  ( .D(n4767), .CK(clk), .RN(n538), .Q(
        \CACHE[1][118] ), .QN(n6007) );
  DFFRX1 \CACHE_reg[1][117]  ( .D(n4768), .CK(clk), .RN(n539), .Q(
        \CACHE[1][117] ), .QN(n6008) );
  DFFRX1 \CACHE_reg[1][116]  ( .D(n4769), .CK(clk), .RN(n540), .Q(
        \CACHE[1][116] ), .QN(n6009) );
  DFFRX1 \CACHE_reg[1][115]  ( .D(n4770), .CK(clk), .RN(n540), .Q(
        \CACHE[1][115] ), .QN(n6010) );
  DFFRX1 \CACHE_reg[1][114]  ( .D(n4771), .CK(clk), .RN(n3020), .Q(
        \CACHE[1][114] ), .QN(n6011) );
  DFFRX1 \CACHE_reg[1][113]  ( .D(n4772), .CK(clk), .RN(n3022), .Q(
        \CACHE[1][113] ), .QN(n6012) );
  DFFRX1 \CACHE_reg[1][112]  ( .D(n4773), .CK(clk), .RN(n3022), .Q(
        \CACHE[1][112] ), .QN(n6013) );
  DFFRX1 \CACHE_reg[1][111]  ( .D(n4774), .CK(clk), .RN(n3023), .Q(
        \CACHE[1][111] ), .QN(n6014) );
  DFFRX1 \CACHE_reg[1][110]  ( .D(n4775), .CK(clk), .RN(n3024), .Q(
        \CACHE[1][110] ), .QN(n6015) );
  DFFRX1 \CACHE_reg[1][109]  ( .D(n4776), .CK(clk), .RN(n3024), .Q(
        \CACHE[1][109] ), .QN(n6016) );
  DFFRX1 \CACHE_reg[1][108]  ( .D(n4777), .CK(clk), .RN(n3025), .Q(
        \CACHE[1][108] ), .QN(n6017) );
  DFFRX1 \CACHE_reg[1][107]  ( .D(n4778), .CK(clk), .RN(n3026), .Q(
        \CACHE[1][107] ), .QN(n6018) );
  DFFRX1 \CACHE_reg[1][106]  ( .D(n4779), .CK(clk), .RN(n3026), .Q(
        \CACHE[1][106] ), .QN(n6019) );
  DFFRX1 \CACHE_reg[1][105]  ( .D(n4780), .CK(clk), .RN(n3027), .Q(
        \CACHE[1][105] ), .QN(n6020) );
  DFFRX1 \CACHE_reg[1][104]  ( .D(n4781), .CK(clk), .RN(n3028), .Q(
        \CACHE[1][104] ), .QN(n6021) );
  DFFRX1 \CACHE_reg[1][103]  ( .D(n4782), .CK(clk), .RN(n3028), .Q(
        \CACHE[1][103] ), .QN(n6022) );
  DFFRX1 \CACHE_reg[1][102]  ( .D(n4783), .CK(clk), .RN(n3029), .Q(
        \CACHE[1][102] ), .QN(n6023) );
  DFFRX1 \CACHE_reg[1][101]  ( .D(n4784), .CK(clk), .RN(n3030), .Q(
        \CACHE[1][101] ), .QN(n6024) );
  DFFRX1 \CACHE_reg[1][100]  ( .D(n4785), .CK(clk), .RN(n3030), .Q(
        \CACHE[1][100] ), .QN(n6025) );
  DFFRX1 \CACHE_reg[1][99]  ( .D(n4786), .CK(clk), .RN(n3031), .Q(
        \CACHE[1][99] ), .QN(n6026) );
  DFFRX1 \CACHE_reg[1][98]  ( .D(n4787), .CK(clk), .RN(n3032), .Q(
        \CACHE[1][98] ), .QN(n6027) );
  DFFRX1 \CACHE_reg[1][97]  ( .D(n4788), .CK(clk), .RN(n3032), .Q(
        \CACHE[1][97] ), .QN(n6028) );
  DFFRX1 \CACHE_reg[1][96]  ( .D(n4789), .CK(clk), .RN(n3033), .Q(
        \CACHE[1][96] ), .QN(n6029) );
  DFFRX1 \CACHE_reg[1][95]  ( .D(n4790), .CK(clk), .RN(n3034), .Q(
        \CACHE[1][95] ), .QN(n6030) );
  DFFRX1 \CACHE_reg[1][94]  ( .D(n4791), .CK(clk), .RN(n3034), .Q(
        \CACHE[1][94] ), .QN(n6031) );
  DFFRX1 \CACHE_reg[1][93]  ( .D(n4792), .CK(clk), .RN(n3035), .Q(
        \CACHE[1][93] ), .QN(n6032) );
  DFFRX1 \CACHE_reg[1][92]  ( .D(n4793), .CK(clk), .RN(n3036), .Q(
        \CACHE[1][92] ), .QN(n6033) );
  DFFRX1 \CACHE_reg[1][91]  ( .D(n4794), .CK(clk), .RN(n3036), .Q(
        \CACHE[1][91] ), .QN(n6034) );
  DFFRX1 \CACHE_reg[1][90]  ( .D(n4795), .CK(clk), .RN(n3037), .Q(
        \CACHE[1][90] ), .QN(n6035) );
  DFFRX1 \CACHE_reg[1][89]  ( .D(n4796), .CK(clk), .RN(n3038), .Q(
        \CACHE[1][89] ), .QN(n6036) );
  DFFRX1 \CACHE_reg[1][88]  ( .D(n4797), .CK(clk), .RN(n3038), .Q(
        \CACHE[1][88] ), .QN(n6037) );
  DFFRX1 \CACHE_reg[1][87]  ( .D(n4798), .CK(clk), .RN(n3039), .Q(
        \CACHE[1][87] ), .QN(n6038) );
  DFFRX1 \CACHE_reg[1][86]  ( .D(n4799), .CK(clk), .RN(n3040), .Q(
        \CACHE[1][86] ), .QN(n6039) );
  DFFRX1 \CACHE_reg[1][85]  ( .D(n4800), .CK(clk), .RN(n3040), .Q(
        \CACHE[1][85] ), .QN(n6040) );
  DFFRX1 \CACHE_reg[1][84]  ( .D(n4801), .CK(clk), .RN(n3041), .Q(
        \CACHE[1][84] ), .QN(n6041) );
  DFFRX1 \CACHE_reg[1][83]  ( .D(n4802), .CK(clk), .RN(n3042), .Q(
        \CACHE[1][83] ), .QN(n6042) );
  DFFRX1 \CACHE_reg[1][82]  ( .D(n4803), .CK(clk), .RN(n3042), .Q(
        \CACHE[1][82] ), .QN(n6043) );
  DFFRX1 \CACHE_reg[1][81]  ( .D(n4804), .CK(clk), .RN(n3043), .Q(
        \CACHE[1][81] ), .QN(n6044) );
  DFFRX1 \CACHE_reg[1][80]  ( .D(n4805), .CK(clk), .RN(n3044), .Q(
        \CACHE[1][80] ), .QN(n6045) );
  DFFRX1 \CACHE_reg[1][79]  ( .D(n4806), .CK(clk), .RN(n3044), .Q(
        \CACHE[1][79] ), .QN(n6046) );
  DFFRX1 \CACHE_reg[1][78]  ( .D(n4807), .CK(clk), .RN(n3045), .Q(
        \CACHE[1][78] ), .QN(n6047) );
  DFFRX1 \CACHE_reg[1][77]  ( .D(n4808), .CK(clk), .RN(n3046), .Q(
        \CACHE[1][77] ), .QN(n6048) );
  DFFRX1 \CACHE_reg[1][76]  ( .D(n4809), .CK(clk), .RN(n3046), .Q(
        \CACHE[1][76] ), .QN(n6049) );
  DFFRX1 \CACHE_reg[1][75]  ( .D(n4810), .CK(clk), .RN(n3047), .Q(
        \CACHE[1][75] ), .QN(n6050) );
  DFFRX1 \CACHE_reg[1][74]  ( .D(n4811), .CK(clk), .RN(n3048), .Q(
        \CACHE[1][74] ), .QN(n6051) );
  DFFRX1 \CACHE_reg[1][73]  ( .D(n4812), .CK(clk), .RN(n3048), .Q(
        \CACHE[1][73] ), .QN(n6052) );
  DFFRX1 \CACHE_reg[1][72]  ( .D(n4813), .CK(clk), .RN(n3049), .Q(
        \CACHE[1][72] ), .QN(n6053) );
  DFFRX1 \CACHE_reg[1][71]  ( .D(n4814), .CK(clk), .RN(n3050), .Q(
        \CACHE[1][71] ), .QN(n6054) );
  DFFRX1 \CACHE_reg[1][70]  ( .D(n4815), .CK(clk), .RN(n3050), .Q(
        \CACHE[1][70] ), .QN(n6055) );
  DFFRX1 \CACHE_reg[1][69]  ( .D(n4816), .CK(clk), .RN(n3051), .Q(
        \CACHE[1][69] ), .QN(n6056) );
  DFFRX1 \CACHE_reg[1][68]  ( .D(n4817), .CK(clk), .RN(n3052), .Q(
        \CACHE[1][68] ), .QN(n6057) );
  DFFRX1 \CACHE_reg[1][67]  ( .D(n4818), .CK(clk), .RN(n3052), .Q(
        \CACHE[1][67] ), .QN(n6058) );
  DFFRX1 \CACHE_reg[1][66]  ( .D(n4819), .CK(clk), .RN(n3053), .Q(
        \CACHE[1][66] ), .QN(n6059) );
  DFFRX1 \CACHE_reg[1][65]  ( .D(n4820), .CK(clk), .RN(n3054), .Q(
        \CACHE[1][65] ), .QN(n6060) );
  DFFRX1 \CACHE_reg[1][64]  ( .D(n4821), .CK(clk), .RN(n3054), .Q(
        \CACHE[1][64] ), .QN(n6061) );
  DFFRX1 \CACHE_reg[1][63]  ( .D(n4822), .CK(clk), .RN(n513), .Q(
        \CACHE[1][63] ), .QN(n6062) );
  DFFRX1 \CACHE_reg[1][62]  ( .D(n4823), .CK(clk), .RN(n513), .Q(
        \CACHE[1][62] ), .QN(n6063) );
  DFFRX1 \CACHE_reg[1][61]  ( .D(n4824), .CK(clk), .RN(n514), .Q(
        \CACHE[1][61] ), .QN(n6064) );
  DFFRX1 \CACHE_reg[1][60]  ( .D(n4825), .CK(clk), .RN(n515), .Q(
        \CACHE[1][60] ), .QN(n6065) );
  DFFRX1 \CACHE_reg[1][59]  ( .D(n4826), .CK(clk), .RN(n515), .Q(
        \CACHE[1][59] ), .QN(n6066) );
  DFFRX1 \CACHE_reg[1][58]  ( .D(n4827), .CK(clk), .RN(n516), .Q(
        \CACHE[1][58] ), .QN(n6067) );
  DFFRX1 \CACHE_reg[1][57]  ( .D(n4828), .CK(clk), .RN(n517), .Q(
        \CACHE[1][57] ), .QN(n6068) );
  DFFRX1 \CACHE_reg[1][56]  ( .D(n4829), .CK(clk), .RN(n517), .Q(
        \CACHE[1][56] ), .QN(n6069) );
  DFFRX1 \CACHE_reg[1][55]  ( .D(n4830), .CK(clk), .RN(n518), .Q(
        \CACHE[1][55] ), .QN(n6070) );
  DFFRX1 \CACHE_reg[1][54]  ( .D(n4831), .CK(clk), .RN(n519), .Q(
        \CACHE[1][54] ), .QN(n6071) );
  DFFRX1 \CACHE_reg[1][53]  ( .D(n4832), .CK(clk), .RN(n519), .Q(
        \CACHE[1][53] ), .QN(n6072) );
  DFFRX1 \CACHE_reg[1][52]  ( .D(n4833), .CK(clk), .RN(n520), .Q(
        \CACHE[1][52] ), .QN(n6073) );
  DFFRX1 \CACHE_reg[1][51]  ( .D(n4834), .CK(clk), .RN(n521), .Q(
        \CACHE[1][51] ), .QN(n6074) );
  DFFRX1 \CACHE_reg[1][50]  ( .D(n4835), .CK(clk), .RN(n521), .Q(
        \CACHE[1][50] ), .QN(n6075) );
  DFFRX1 \CACHE_reg[1][49]  ( .D(n4836), .CK(clk), .RN(n522), .Q(
        \CACHE[1][49] ), .QN(n6076) );
  DFFRX1 \CACHE_reg[1][48]  ( .D(n4837), .CK(clk), .RN(n523), .Q(
        \CACHE[1][48] ), .QN(n6077) );
  DFFRX1 \CACHE_reg[1][47]  ( .D(n4838), .CK(clk), .RN(n523), .Q(
        \CACHE[1][47] ), .QN(n6078) );
  DFFRX1 \CACHE_reg[1][46]  ( .D(n4839), .CK(clk), .RN(n524), .Q(
        \CACHE[1][46] ), .QN(n6079) );
  DFFRX1 \CACHE_reg[1][45]  ( .D(n4840), .CK(clk), .RN(n525), .Q(
        \CACHE[1][45] ), .QN(n6080) );
  DFFRX1 \CACHE_reg[1][44]  ( .D(n4841), .CK(clk), .RN(n525), .Q(
        \CACHE[1][44] ), .QN(n6081) );
  DFFRX1 \CACHE_reg[1][43]  ( .D(n4842), .CK(clk), .RN(n526), .Q(
        \CACHE[1][43] ), .QN(n6082) );
  DFFRX1 \CACHE_reg[1][42]  ( .D(n4843), .CK(clk), .RN(n527), .Q(
        \CACHE[1][42] ), .QN(n6083) );
  DFFRX1 \CACHE_reg[1][41]  ( .D(n4844), .CK(clk), .RN(n527), .Q(
        \CACHE[1][41] ), .QN(n6084) );
  DFFRX1 \CACHE_reg[1][40]  ( .D(n4845), .CK(clk), .RN(n528), .Q(
        \CACHE[1][40] ), .QN(n6085) );
  DFFRX1 \CACHE_reg[1][39]  ( .D(n4846), .CK(clk), .RN(n529), .Q(
        \CACHE[1][39] ), .QN(n6086) );
  DFFRX1 \CACHE_reg[1][38]  ( .D(n4847), .CK(clk), .RN(n529), .Q(
        \CACHE[1][38] ), .QN(n6087) );
  DFFRX1 \CACHE_reg[1][37]  ( .D(n4848), .CK(clk), .RN(n530), .Q(
        \CACHE[1][37] ), .QN(n6088) );
  DFFRX1 \CACHE_reg[1][36]  ( .D(n4849), .CK(clk), .RN(n531), .Q(
        \CACHE[1][36] ), .QN(n6089) );
  DFFRX1 \CACHE_reg[1][35]  ( .D(n4850), .CK(clk), .RN(n531), .Q(
        \CACHE[1][35] ), .QN(n6090) );
  DFFRX1 \CACHE_reg[1][34]  ( .D(n4851), .CK(clk), .RN(n532), .Q(
        \CACHE[1][34] ), .QN(n6091) );
  DFFRX1 \CACHE_reg[1][33]  ( .D(n4852), .CK(clk), .RN(n533), .Q(
        \CACHE[1][33] ), .QN(n6092) );
  DFFRX1 \CACHE_reg[1][32]  ( .D(n4853), .CK(clk), .RN(n533), .Q(
        \CACHE[1][32] ), .QN(n6093) );
  DFFRX1 \CACHE_reg[1][31]  ( .D(n4854), .CK(clk), .RN(n491), .Q(
        \CACHE[1][31] ), .QN(n6094) );
  DFFRX1 \CACHE_reg[1][30]  ( .D(n4855), .CK(clk), .RN(n3055), .Q(
        \CACHE[1][30] ), .QN(n6095) );
  DFFRX1 \CACHE_reg[1][29]  ( .D(n4856), .CK(clk), .RN(n493), .Q(
        \CACHE[1][29] ), .QN(n6096) );
  DFFRX1 \CACHE_reg[1][28]  ( .D(n4857), .CK(clk), .RN(n493), .Q(
        \CACHE[1][28] ), .QN(n6097) );
  DFFRX1 \CACHE_reg[1][27]  ( .D(n4858), .CK(clk), .RN(n494), .Q(
        \CACHE[1][27] ), .QN(n6098) );
  DFFRX1 \CACHE_reg[1][26]  ( .D(n4859), .CK(clk), .RN(n495), .Q(
        \CACHE[1][26] ), .QN(n6099) );
  DFFRX1 \CACHE_reg[1][25]  ( .D(n4860), .CK(clk), .RN(n495), .Q(
        \CACHE[1][25] ), .QN(n6100) );
  DFFRX1 \CACHE_reg[1][24]  ( .D(n4861), .CK(clk), .RN(n496), .Q(
        \CACHE[1][24] ), .QN(n6101) );
  DFFRX1 \CACHE_reg[1][23]  ( .D(n4862), .CK(clk), .RN(n497), .Q(
        \CACHE[1][23] ), .QN(n6102) );
  DFFRX1 \CACHE_reg[1][22]  ( .D(n4863), .CK(clk), .RN(n497), .Q(
        \CACHE[1][22] ), .QN(n6103) );
  DFFRX1 \CACHE_reg[1][21]  ( .D(n4864), .CK(clk), .RN(n498), .Q(
        \CACHE[1][21] ), .QN(n6104) );
  DFFRX1 \CACHE_reg[1][20]  ( .D(n4865), .CK(clk), .RN(n499), .Q(
        \CACHE[1][20] ), .QN(n6105) );
  DFFRX1 \CACHE_reg[1][19]  ( .D(n4866), .CK(clk), .RN(n499), .Q(
        \CACHE[1][19] ), .QN(n6106) );
  DFFRX1 \CACHE_reg[1][18]  ( .D(n4867), .CK(clk), .RN(n500), .Q(
        \CACHE[1][18] ), .QN(n6107) );
  DFFRX1 \CACHE_reg[1][17]  ( .D(n4868), .CK(clk), .RN(n501), .Q(
        \CACHE[1][17] ), .QN(n6108) );
  DFFRX1 \CACHE_reg[1][16]  ( .D(n4869), .CK(clk), .RN(n501), .Q(
        \CACHE[1][16] ), .QN(n6109) );
  DFFRX1 \CACHE_reg[1][15]  ( .D(n4870), .CK(clk), .RN(n502), .Q(
        \CACHE[1][15] ), .QN(n6110) );
  DFFRX1 \CACHE_reg[1][14]  ( .D(n4871), .CK(clk), .RN(n503), .Q(
        \CACHE[1][14] ), .QN(n6111) );
  DFFRX1 \CACHE_reg[1][13]  ( .D(n4872), .CK(clk), .RN(n503), .Q(
        \CACHE[1][13] ), .QN(n6112) );
  DFFRX1 \CACHE_reg[1][12]  ( .D(n4873), .CK(clk), .RN(n504), .Q(
        \CACHE[1][12] ), .QN(n6113) );
  DFFRX1 \CACHE_reg[1][11]  ( .D(n4874), .CK(clk), .RN(n505), .Q(
        \CACHE[1][11] ), .QN(n6114) );
  DFFRX1 \CACHE_reg[1][10]  ( .D(n4875), .CK(clk), .RN(n505), .Q(
        \CACHE[1][10] ), .QN(n6115) );
  DFFRX1 \CACHE_reg[1][9]  ( .D(n4876), .CK(clk), .RN(n506), .Q(\CACHE[1][9] ), 
        .QN(n6116) );
  DFFRX1 \CACHE_reg[1][8]  ( .D(n4877), .CK(clk), .RN(n507), .Q(\CACHE[1][8] ), 
        .QN(n6117) );
  DFFRX1 \CACHE_reg[1][7]  ( .D(n4878), .CK(clk), .RN(n507), .Q(\CACHE[1][7] ), 
        .QN(n6118) );
  DFFRX1 \CACHE_reg[1][6]  ( .D(n4879), .CK(clk), .RN(n508), .Q(\CACHE[1][6] ), 
        .QN(n6119) );
  DFFRX1 \CACHE_reg[1][5]  ( .D(n4880), .CK(clk), .RN(n509), .Q(\CACHE[1][5] ), 
        .QN(n6120) );
  DFFRX1 \CACHE_reg[1][4]  ( .D(n4881), .CK(clk), .RN(n509), .Q(\CACHE[1][4] ), 
        .QN(n6121) );
  DFFRX1 \CACHE_reg[1][3]  ( .D(n4882), .CK(clk), .RN(n510), .Q(\CACHE[1][3] ), 
        .QN(n6122) );
  DFFRX1 \CACHE_reg[1][2]  ( .D(n4883), .CK(clk), .RN(n511), .Q(\CACHE[1][2] ), 
        .QN(n6123) );
  DFFRX1 \CACHE_reg[1][1]  ( .D(n4884), .CK(clk), .RN(n511), .Q(\CACHE[1][1] ), 
        .QN(n6124) );
  DFFRX1 \CACHE_reg[1][0]  ( .D(n4885), .CK(clk), .RN(n512), .Q(\CACHE[1][0] ), 
        .QN(n6125) );
  DFFRX1 \CACHE_reg[4][154]  ( .D(n4266), .CK(clk), .RN(n3056), .Q(
        \CACHE[4][154] ), .QN(n5506) );
  DFFRX1 \CACHE_reg[4][153]  ( .D(n4267), .CK(clk), .RN(n3056), .Q(
        \CACHE[4][153] ), .QN(n5507) );
  DFFRX1 \CACHE_reg[4][152]  ( .D(n4268), .CK(clk), .RN(n474), .Q(
        \CACHE[4][152] ), .QN(n5508) );
  DFFRX1 \CACHE_reg[4][151]  ( .D(n4269), .CK(clk), .RN(n475), .Q(
        \CACHE[4][151] ), .QN(n5509) );
  DFFRX1 \CACHE_reg[4][150]  ( .D(n4270), .CK(clk), .RN(n476), .Q(
        \CACHE[4][150] ), .QN(n5510) );
  DFFRX1 \CACHE_reg[4][149]  ( .D(n4271), .CK(clk), .RN(n476), .Q(
        \CACHE[4][149] ), .QN(n5511) );
  DFFRX1 \CACHE_reg[4][148]  ( .D(n4272), .CK(clk), .RN(n477), .Q(
        \CACHE[4][148] ), .QN(n5512) );
  DFFRX1 \CACHE_reg[4][147]  ( .D(n4273), .CK(clk), .RN(n478), .Q(
        \CACHE[4][147] ), .QN(n5513) );
  DFFRX1 \CACHE_reg[4][146]  ( .D(n4274), .CK(clk), .RN(n478), .Q(
        \CACHE[4][146] ), .QN(n5514) );
  DFFRX1 \CACHE_reg[4][145]  ( .D(n4275), .CK(clk), .RN(n479), .Q(
        \CACHE[4][145] ), .QN(n5515) );
  DFFRX1 \CACHE_reg[4][144]  ( .D(n4276), .CK(clk), .RN(n480), .Q(
        \CACHE[4][144] ), .QN(n5516) );
  DFFRX1 \CACHE_reg[4][143]  ( .D(n4277), .CK(clk), .RN(n480), .Q(
        \CACHE[4][143] ), .QN(n5517) );
  DFFRX1 \CACHE_reg[4][142]  ( .D(n4278), .CK(clk), .RN(n481), .Q(
        \CACHE[4][142] ), .QN(n5518) );
  DFFRX1 \CACHE_reg[4][141]  ( .D(n4279), .CK(clk), .RN(n482), .Q(
        \CACHE[4][141] ), .QN(n5519) );
  DFFRX1 \CACHE_reg[4][140]  ( .D(n4280), .CK(clk), .RN(n482), .Q(
        \CACHE[4][140] ), .QN(n5520) );
  DFFRX1 \CACHE_reg[4][139]  ( .D(n4281), .CK(clk), .RN(n490), .Q(
        \CACHE[4][139] ), .QN(n5521) );
  DFFRX1 \CACHE_reg[4][138]  ( .D(n4282), .CK(clk), .RN(n483), .Q(
        \CACHE[4][138] ), .QN(n5522) );
  DFFRX1 \CACHE_reg[4][137]  ( .D(n4283), .CK(clk), .RN(n484), .Q(
        \CACHE[4][137] ), .QN(n5523) );
  DFFRX1 \CACHE_reg[4][136]  ( .D(n4284), .CK(clk), .RN(n484), .Q(
        \CACHE[4][136] ), .QN(n5524) );
  DFFRX1 \CACHE_reg[4][135]  ( .D(n4285), .CK(clk), .RN(n485), .Q(
        \CACHE[4][135] ), .QN(n5525) );
  DFFRX1 \CACHE_reg[4][134]  ( .D(n4286), .CK(clk), .RN(n486), .Q(
        \CACHE[4][134] ), .QN(n5526) );
  DFFRX1 \CACHE_reg[4][133]  ( .D(n4287), .CK(clk), .RN(n486), .Q(
        \CACHE[4][133] ), .QN(n5527) );
  DFFRX1 \CACHE_reg[4][132]  ( .D(n4288), .CK(clk), .RN(n474), .Q(
        \CACHE[4][132] ), .QN(n5528) );
  DFFRX1 \CACHE_reg[4][131]  ( .D(n4289), .CK(clk), .RN(n487), .Q(
        \CACHE[4][131] ), .QN(n5529) );
  DFFRX1 \CACHE_reg[4][130]  ( .D(n4290), .CK(clk), .RN(n488), .Q(
        \CACHE[4][130] ), .QN(n5530) );
  DFFRX1 \CACHE_reg[4][129]  ( .D(n4291), .CK(clk), .RN(n488), .Q(
        \CACHE[4][129] ), .QN(n5531) );
  DFFRX1 \CACHE_reg[4][128]  ( .D(n4292), .CK(clk), .RN(n489), .Q(
        \CACHE[4][128] ), .QN(n5532) );
  DFFRX1 \CACHE_reg[4][127]  ( .D(n4293), .CK(clk), .RN(n3056), .Q(
        \CACHE[4][127] ), .QN(n5533) );
  DFFRX1 \CACHE_reg[4][126]  ( .D(n4294), .CK(clk), .RN(n491), .Q(
        \CACHE[4][126] ), .QN(n5534) );
  DFFRX1 \CACHE_reg[4][125]  ( .D(n4295), .CK(clk), .RN(n534), .Q(
        \CACHE[4][125] ), .QN(n5535) );
  DFFRX1 \CACHE_reg[4][124]  ( .D(n4296), .CK(clk), .RN(n534), .Q(
        \CACHE[4][124] ), .QN(n5536) );
  DFFRX1 \CACHE_reg[4][123]  ( .D(n4297), .CK(clk), .RN(n535), .Q(
        \CACHE[4][123] ), .QN(n5537) );
  DFFRX1 \CACHE_reg[4][122]  ( .D(n4298), .CK(clk), .RN(n535), .Q(
        \CACHE[4][122] ), .QN(n5538) );
  DFFRX1 \CACHE_reg[4][121]  ( .D(n4299), .CK(clk), .RN(n536), .Q(
        \CACHE[4][121] ), .QN(n5539) );
  DFFRX1 \CACHE_reg[4][120]  ( .D(n4300), .CK(clk), .RN(n537), .Q(
        \CACHE[4][120] ), .QN(n5540) );
  DFFRX1 \CACHE_reg[4][119]  ( .D(n4301), .CK(clk), .RN(n537), .Q(
        \CACHE[4][119] ), .QN(n5541) );
  DFFRX1 \CACHE_reg[4][118]  ( .D(n4302), .CK(clk), .RN(n538), .Q(
        \CACHE[4][118] ), .QN(n5542) );
  DFFRX1 \CACHE_reg[4][117]  ( .D(n4303), .CK(clk), .RN(n539), .Q(
        \CACHE[4][117] ), .QN(n5543) );
  DFFRX1 \CACHE_reg[4][116]  ( .D(n4304), .CK(clk), .RN(n539), .Q(
        \CACHE[4][116] ), .QN(n5544) );
  DFFRX1 \CACHE_reg[4][115]  ( .D(n4305), .CK(clk), .RN(n540), .Q(
        \CACHE[4][115] ), .QN(n5545) );
  DFFRX1 \CACHE_reg[4][114]  ( .D(n4306), .CK(clk), .RN(n3020), .Q(
        \CACHE[4][114] ), .QN(n5546) );
  DFFRX1 \CACHE_reg[4][113]  ( .D(n4307), .CK(clk), .RN(n3020), .Q(
        \CACHE[4][113] ), .QN(n5547) );
  DFFRX1 \CACHE_reg[4][112]  ( .D(n4308), .CK(clk), .RN(n3022), .Q(
        \CACHE[4][112] ), .QN(n5548) );
  DFFRX1 \CACHE_reg[4][111]  ( .D(n4309), .CK(clk), .RN(n3023), .Q(
        \CACHE[4][111] ), .QN(n5549) );
  DFFRX1 \CACHE_reg[4][110]  ( .D(n4310), .CK(clk), .RN(n3023), .Q(
        \CACHE[4][110] ), .QN(n5550) );
  DFFRX1 \CACHE_reg[4][109]  ( .D(n4311), .CK(clk), .RN(n3024), .Q(
        \CACHE[4][109] ), .QN(n5551) );
  DFFRX1 \CACHE_reg[4][108]  ( .D(n4312), .CK(clk), .RN(n3025), .Q(
        \CACHE[4][108] ), .QN(n5552) );
  DFFRX1 \CACHE_reg[4][107]  ( .D(n4313), .CK(clk), .RN(n3025), .Q(
        \CACHE[4][107] ), .QN(n5553) );
  DFFRX1 \CACHE_reg[4][106]  ( .D(n4314), .CK(clk), .RN(n3026), .Q(
        \CACHE[4][106] ), .QN(n5554) );
  DFFRX1 \CACHE_reg[4][105]  ( .D(n4315), .CK(clk), .RN(n3027), .Q(
        \CACHE[4][105] ), .QN(n5555) );
  DFFRX1 \CACHE_reg[4][104]  ( .D(n4316), .CK(clk), .RN(n3027), .Q(
        \CACHE[4][104] ), .QN(n5556) );
  DFFRX1 \CACHE_reg[4][103]  ( .D(n4317), .CK(clk), .RN(n3028), .Q(
        \CACHE[4][103] ), .QN(n5557) );
  DFFRX1 \CACHE_reg[4][102]  ( .D(n4318), .CK(clk), .RN(n3029), .Q(
        \CACHE[4][102] ), .QN(n5558) );
  DFFRX1 \CACHE_reg[4][101]  ( .D(n4319), .CK(clk), .RN(n3029), .Q(
        \CACHE[4][101] ), .QN(n5559) );
  DFFRX1 \CACHE_reg[4][100]  ( .D(n4320), .CK(clk), .RN(n3030), .Q(
        \CACHE[4][100] ), .QN(n5560) );
  DFFRX1 \CACHE_reg[4][99]  ( .D(n4321), .CK(clk), .RN(n3031), .Q(
        \CACHE[4][99] ), .QN(n5561) );
  DFFRX1 \CACHE_reg[4][98]  ( .D(n4322), .CK(clk), .RN(n3031), .Q(
        \CACHE[4][98] ), .QN(n5562) );
  DFFRX1 \CACHE_reg[4][97]  ( .D(n4323), .CK(clk), .RN(n3032), .Q(
        \CACHE[4][97] ), .QN(n5563) );
  DFFRX1 \CACHE_reg[4][96]  ( .D(n4324), .CK(clk), .RN(n3033), .Q(
        \CACHE[4][96] ), .QN(n5564) );
  DFFRX1 \CACHE_reg[4][95]  ( .D(n4325), .CK(clk), .RN(n3033), .Q(
        \CACHE[4][95] ), .QN(n5565) );
  DFFRX1 \CACHE_reg[4][94]  ( .D(n4326), .CK(clk), .RN(n3034), .Q(
        \CACHE[4][94] ), .QN(n5566) );
  DFFRX1 \CACHE_reg[4][93]  ( .D(n4327), .CK(clk), .RN(n3035), .Q(
        \CACHE[4][93] ), .QN(n5567) );
  DFFRX1 \CACHE_reg[4][92]  ( .D(n4328), .CK(clk), .RN(n3035), .Q(
        \CACHE[4][92] ), .QN(n5568) );
  DFFRX1 \CACHE_reg[4][91]  ( .D(n4329), .CK(clk), .RN(n3036), .Q(
        \CACHE[4][91] ), .QN(n5569) );
  DFFRX1 \CACHE_reg[4][90]  ( .D(n4330), .CK(clk), .RN(n3037), .Q(
        \CACHE[4][90] ), .QN(n5570) );
  DFFRX1 \CACHE_reg[4][89]  ( .D(n4331), .CK(clk), .RN(n3037), .Q(
        \CACHE[4][89] ), .QN(n5571) );
  DFFRX1 \CACHE_reg[4][88]  ( .D(n4332), .CK(clk), .RN(n3038), .Q(
        \CACHE[4][88] ), .QN(n5572) );
  DFFRX1 \CACHE_reg[4][87]  ( .D(n4333), .CK(clk), .RN(n3039), .Q(
        \CACHE[4][87] ), .QN(n5573) );
  DFFRX1 \CACHE_reg[4][86]  ( .D(n4334), .CK(clk), .RN(n3039), .Q(
        \CACHE[4][86] ), .QN(n5574) );
  DFFRX1 \CACHE_reg[4][85]  ( .D(n4335), .CK(clk), .RN(n3040), .Q(
        \CACHE[4][85] ), .QN(n5575) );
  DFFRX1 \CACHE_reg[4][84]  ( .D(n4336), .CK(clk), .RN(n3041), .Q(
        \CACHE[4][84] ), .QN(n5576) );
  DFFRX1 \CACHE_reg[4][83]  ( .D(n4337), .CK(clk), .RN(n3041), .Q(
        \CACHE[4][83] ), .QN(n5577) );
  DFFRX1 \CACHE_reg[4][82]  ( .D(n4338), .CK(clk), .RN(n3042), .Q(
        \CACHE[4][82] ), .QN(n5578) );
  DFFRX1 \CACHE_reg[4][81]  ( .D(n4339), .CK(clk), .RN(n3043), .Q(
        \CACHE[4][81] ), .QN(n5579) );
  DFFRX1 \CACHE_reg[4][80]  ( .D(n4340), .CK(clk), .RN(n3043), .Q(
        \CACHE[4][80] ), .QN(n5580) );
  DFFRX1 \CACHE_reg[4][79]  ( .D(n4341), .CK(clk), .RN(n3044), .Q(
        \CACHE[4][79] ), .QN(n5581) );
  DFFRX1 \CACHE_reg[4][78]  ( .D(n4342), .CK(clk), .RN(n3045), .Q(
        \CACHE[4][78] ), .QN(n5582) );
  DFFRX1 \CACHE_reg[4][77]  ( .D(n4343), .CK(clk), .RN(n3045), .Q(
        \CACHE[4][77] ), .QN(n5583) );
  DFFRX1 \CACHE_reg[4][76]  ( .D(n4344), .CK(clk), .RN(n3046), .Q(
        \CACHE[4][76] ), .QN(n5584) );
  DFFRX1 \CACHE_reg[4][75]  ( .D(n4345), .CK(clk), .RN(n3047), .Q(
        \CACHE[4][75] ), .QN(n5585) );
  DFFRX1 \CACHE_reg[4][74]  ( .D(n4346), .CK(clk), .RN(n3047), .Q(
        \CACHE[4][74] ), .QN(n5586) );
  DFFRX1 \CACHE_reg[4][73]  ( .D(n4347), .CK(clk), .RN(n3048), .Q(
        \CACHE[4][73] ), .QN(n5587) );
  DFFRX1 \CACHE_reg[4][72]  ( .D(n4348), .CK(clk), .RN(n3049), .Q(
        \CACHE[4][72] ), .QN(n5588) );
  DFFRX1 \CACHE_reg[4][71]  ( .D(n4349), .CK(clk), .RN(n3049), .Q(
        \CACHE[4][71] ), .QN(n5589) );
  DFFRX1 \CACHE_reg[4][70]  ( .D(n4350), .CK(clk), .RN(n3050), .Q(
        \CACHE[4][70] ), .QN(n5590) );
  DFFRX1 \CACHE_reg[4][69]  ( .D(n4351), .CK(clk), .RN(n3051), .Q(
        \CACHE[4][69] ), .QN(n5591) );
  DFFRX1 \CACHE_reg[4][68]  ( .D(n4352), .CK(clk), .RN(n3051), .Q(
        \CACHE[4][68] ), .QN(n5592) );
  DFFRX1 \CACHE_reg[4][67]  ( .D(n4353), .CK(clk), .RN(n3052), .Q(
        \CACHE[4][67] ), .QN(n5593) );
  DFFRX1 \CACHE_reg[4][66]  ( .D(n4354), .CK(clk), .RN(n3053), .Q(
        \CACHE[4][66] ), .QN(n5594) );
  DFFRX1 \CACHE_reg[4][65]  ( .D(n4355), .CK(clk), .RN(n3053), .Q(
        \CACHE[4][65] ), .QN(n5595) );
  DFFRX1 \CACHE_reg[4][64]  ( .D(n4356), .CK(clk), .RN(n3054), .Q(
        \CACHE[4][64] ), .QN(n5596) );
  DFFRX1 \CACHE_reg[4][63]  ( .D(n4357), .CK(clk), .RN(n512), .Q(
        \CACHE[4][63] ), .QN(n5597) );
  DFFRX1 \CACHE_reg[4][62]  ( .D(n4358), .CK(clk), .RN(n513), .Q(
        \CACHE[4][62] ), .QN(n5598) );
  DFFRX1 \CACHE_reg[4][61]  ( .D(n4359), .CK(clk), .RN(n514), .Q(
        \CACHE[4][61] ), .QN(n5599) );
  DFFRX1 \CACHE_reg[4][60]  ( .D(n4360), .CK(clk), .RN(n514), .Q(
        \CACHE[4][60] ), .QN(n5600) );
  DFFRX1 \CACHE_reg[4][59]  ( .D(n4361), .CK(clk), .RN(n515), .Q(
        \CACHE[4][59] ), .QN(n5601) );
  DFFRX1 \CACHE_reg[4][58]  ( .D(n4362), .CK(clk), .RN(n516), .Q(
        \CACHE[4][58] ), .QN(n5602) );
  DFFRX1 \CACHE_reg[4][57]  ( .D(n4363), .CK(clk), .RN(n516), .Q(
        \CACHE[4][57] ), .QN(n5603) );
  DFFRX1 \CACHE_reg[4][56]  ( .D(n4364), .CK(clk), .RN(n517), .Q(
        \CACHE[4][56] ), .QN(n5604) );
  DFFRX1 \CACHE_reg[4][55]  ( .D(n4365), .CK(clk), .RN(n518), .Q(
        \CACHE[4][55] ), .QN(n5605) );
  DFFRX1 \CACHE_reg[4][54]  ( .D(n4366), .CK(clk), .RN(n518), .Q(
        \CACHE[4][54] ), .QN(n5606) );
  DFFRX1 \CACHE_reg[4][53]  ( .D(n4367), .CK(clk), .RN(n519), .Q(
        \CACHE[4][53] ), .QN(n5607) );
  DFFRX1 \CACHE_reg[4][52]  ( .D(n4368), .CK(clk), .RN(n520), .Q(
        \CACHE[4][52] ), .QN(n5608) );
  DFFRX1 \CACHE_reg[4][51]  ( .D(n4369), .CK(clk), .RN(n520), .Q(
        \CACHE[4][51] ), .QN(n5609) );
  DFFRX1 \CACHE_reg[4][50]  ( .D(n4370), .CK(clk), .RN(n521), .Q(
        \CACHE[4][50] ), .QN(n5610) );
  DFFRX1 \CACHE_reg[4][49]  ( .D(n4371), .CK(clk), .RN(n522), .Q(
        \CACHE[4][49] ), .QN(n5611) );
  DFFRX1 \CACHE_reg[4][48]  ( .D(n4372), .CK(clk), .RN(n522), .Q(
        \CACHE[4][48] ), .QN(n5612) );
  DFFRX1 \CACHE_reg[4][47]  ( .D(n4373), .CK(clk), .RN(n523), .Q(
        \CACHE[4][47] ), .QN(n5613) );
  DFFRX1 \CACHE_reg[4][46]  ( .D(n4374), .CK(clk), .RN(n524), .Q(
        \CACHE[4][46] ), .QN(n5614) );
  DFFRX1 \CACHE_reg[4][45]  ( .D(n4375), .CK(clk), .RN(n524), .Q(
        \CACHE[4][45] ), .QN(n5615) );
  DFFRX1 \CACHE_reg[4][44]  ( .D(n4376), .CK(clk), .RN(n525), .Q(
        \CACHE[4][44] ), .QN(n5616) );
  DFFRX1 \CACHE_reg[4][43]  ( .D(n4377), .CK(clk), .RN(n526), .Q(
        \CACHE[4][43] ), .QN(n5617) );
  DFFRX1 \CACHE_reg[4][42]  ( .D(n4378), .CK(clk), .RN(n526), .Q(
        \CACHE[4][42] ), .QN(n5618) );
  DFFRX1 \CACHE_reg[4][41]  ( .D(n4379), .CK(clk), .RN(n527), .Q(
        \CACHE[4][41] ), .QN(n5619) );
  DFFRX1 \CACHE_reg[4][40]  ( .D(n4380), .CK(clk), .RN(n528), .Q(
        \CACHE[4][40] ), .QN(n5620) );
  DFFRX1 \CACHE_reg[4][39]  ( .D(n4381), .CK(clk), .RN(n528), .Q(
        \CACHE[4][39] ), .QN(n5621) );
  DFFRX1 \CACHE_reg[4][38]  ( .D(n4382), .CK(clk), .RN(n529), .Q(
        \CACHE[4][38] ), .QN(n5622) );
  DFFRX1 \CACHE_reg[4][37]  ( .D(n4383), .CK(clk), .RN(n530), .Q(
        \CACHE[4][37] ), .QN(n5623) );
  DFFRX1 \CACHE_reg[4][36]  ( .D(n4384), .CK(clk), .RN(n530), .Q(
        \CACHE[4][36] ), .QN(n5624) );
  DFFRX1 \CACHE_reg[4][35]  ( .D(n4385), .CK(clk), .RN(n531), .Q(
        \CACHE[4][35] ), .QN(n5625) );
  DFFRX1 \CACHE_reg[4][34]  ( .D(n4386), .CK(clk), .RN(n532), .Q(
        \CACHE[4][34] ), .QN(n5626) );
  DFFRX1 \CACHE_reg[4][33]  ( .D(n4387), .CK(clk), .RN(n532), .Q(
        \CACHE[4][33] ), .QN(n5627) );
  DFFRX1 \CACHE_reg[4][32]  ( .D(n4388), .CK(clk), .RN(n533), .Q(
        \CACHE[4][32] ), .QN(n5628) );
  DFFRX1 \CACHE_reg[4][31]  ( .D(n4389), .CK(clk), .RN(n490), .Q(
        \CACHE[4][31] ), .QN(n5629) );
  DFFRX1 \CACHE_reg[4][30]  ( .D(n4390), .CK(clk), .RN(n3056), .Q(
        \CACHE[4][30] ), .QN(n5630) );
  DFFRX1 \CACHE_reg[4][29]  ( .D(n4391), .CK(clk), .RN(n492), .Q(
        \CACHE[4][29] ), .QN(n5631) );
  DFFRX1 \CACHE_reg[4][28]  ( .D(n4392), .CK(clk), .RN(n493), .Q(
        \CACHE[4][28] ), .QN(n5632) );
  DFFRX1 \CACHE_reg[4][27]  ( .D(n4393), .CK(clk), .RN(n494), .Q(
        \CACHE[4][27] ), .QN(n5633) );
  DFFRX1 \CACHE_reg[4][26]  ( .D(n4394), .CK(clk), .RN(n494), .Q(
        \CACHE[4][26] ), .QN(n5634) );
  DFFRX1 \CACHE_reg[4][25]  ( .D(n4395), .CK(clk), .RN(n495), .Q(
        \CACHE[4][25] ), .QN(n5635) );
  DFFRX1 \CACHE_reg[4][24]  ( .D(n4396), .CK(clk), .RN(n496), .Q(
        \CACHE[4][24] ), .QN(n5636) );
  DFFRX1 \CACHE_reg[4][23]  ( .D(n4397), .CK(clk), .RN(n496), .Q(
        \CACHE[4][23] ), .QN(n5637) );
  DFFRX1 \CACHE_reg[4][22]  ( .D(n4398), .CK(clk), .RN(n497), .Q(
        \CACHE[4][22] ), .QN(n5638) );
  DFFRX1 \CACHE_reg[4][21]  ( .D(n4399), .CK(clk), .RN(n498), .Q(
        \CACHE[4][21] ), .QN(n5639) );
  DFFRX1 \CACHE_reg[4][20]  ( .D(n4400), .CK(clk), .RN(n498), .Q(
        \CACHE[4][20] ), .QN(n5640) );
  DFFRX1 \CACHE_reg[4][19]  ( .D(n4401), .CK(clk), .RN(n499), .Q(
        \CACHE[4][19] ), .QN(n5641) );
  DFFRX1 \CACHE_reg[4][18]  ( .D(n4402), .CK(clk), .RN(n500), .Q(
        \CACHE[4][18] ), .QN(n5642) );
  DFFRX1 \CACHE_reg[4][17]  ( .D(n4403), .CK(clk), .RN(n500), .Q(
        \CACHE[4][17] ), .QN(n5643) );
  DFFRX1 \CACHE_reg[4][16]  ( .D(n4404), .CK(clk), .RN(n501), .Q(
        \CACHE[4][16] ), .QN(n5644) );
  DFFRX1 \CACHE_reg[4][15]  ( .D(n4405), .CK(clk), .RN(n502), .Q(
        \CACHE[4][15] ), .QN(n5645) );
  DFFRX1 \CACHE_reg[4][14]  ( .D(n4406), .CK(clk), .RN(n502), .Q(
        \CACHE[4][14] ), .QN(n5646) );
  DFFRX1 \CACHE_reg[4][13]  ( .D(n4407), .CK(clk), .RN(n503), .Q(
        \CACHE[4][13] ), .QN(n5647) );
  DFFRX1 \CACHE_reg[4][12]  ( .D(n4408), .CK(clk), .RN(n504), .Q(
        \CACHE[4][12] ), .QN(n5648) );
  DFFRX1 \CACHE_reg[4][11]  ( .D(n4409), .CK(clk), .RN(n504), .Q(
        \CACHE[4][11] ), .QN(n5649) );
  DFFRX1 \CACHE_reg[4][10]  ( .D(n4410), .CK(clk), .RN(n505), .Q(
        \CACHE[4][10] ), .QN(n5650) );
  DFFRX1 \CACHE_reg[4][9]  ( .D(n4411), .CK(clk), .RN(n506), .Q(\CACHE[4][9] ), 
        .QN(n5651) );
  DFFRX1 \CACHE_reg[4][8]  ( .D(n4412), .CK(clk), .RN(n506), .Q(\CACHE[4][8] ), 
        .QN(n5652) );
  DFFRX1 \CACHE_reg[4][7]  ( .D(n4413), .CK(clk), .RN(n507), .Q(\CACHE[4][7] ), 
        .QN(n5653) );
  DFFRX1 \CACHE_reg[4][6]  ( .D(n4414), .CK(clk), .RN(n508), .Q(\CACHE[4][6] ), 
        .QN(n5654) );
  DFFRX1 \CACHE_reg[4][5]  ( .D(n4415), .CK(clk), .RN(n508), .Q(\CACHE[4][5] ), 
        .QN(n5655) );
  DFFRX1 \CACHE_reg[4][4]  ( .D(n4416), .CK(clk), .RN(n509), .Q(\CACHE[4][4] ), 
        .QN(n5656) );
  DFFRX1 \CACHE_reg[4][3]  ( .D(n4417), .CK(clk), .RN(n510), .Q(\CACHE[4][3] ), 
        .QN(n5657) );
  DFFRX1 \CACHE_reg[4][2]  ( .D(n4418), .CK(clk), .RN(n510), .Q(\CACHE[4][2] ), 
        .QN(n5658) );
  DFFRX1 \CACHE_reg[4][1]  ( .D(n4419), .CK(clk), .RN(n511), .Q(\CACHE[4][1] ), 
        .QN(n5659) );
  DFFRX1 \CACHE_reg[4][0]  ( .D(n4420), .CK(clk), .RN(n512), .Q(\CACHE[4][0] ), 
        .QN(n5660) );
  DFFRX1 \CACHE_reg[0][154]  ( .D(n4886), .CK(clk), .RN(n3055), .Q(
        \CACHE[0][154] ), .QN(n6126) );
  DFFRX1 \CACHE_reg[0][153]  ( .D(n4887), .CK(clk), .RN(n3055), .Q(
        \CACHE[0][153] ), .QN(n6127) );
  DFFRX1 \CACHE_reg[0][152]  ( .D(n4888), .CK(clk), .RN(n475), .Q(
        \CACHE[0][152] ), .QN(n6128) );
  DFFRX1 \CACHE_reg[0][151]  ( .D(n4889), .CK(clk), .RN(n475), .Q(
        \CACHE[0][151] ), .QN(n6129) );
  DFFRX1 \CACHE_reg[0][150]  ( .D(n4890), .CK(clk), .RN(n476), .Q(
        \CACHE[0][150] ), .QN(n6130) );
  DFFRX1 \CACHE_reg[0][149]  ( .D(n4891), .CK(clk), .RN(n477), .Q(
        \CACHE[0][149] ), .QN(n6131) );
  DFFRX1 \CACHE_reg[0][148]  ( .D(n4892), .CK(clk), .RN(n477), .Q(
        \CACHE[0][148] ), .QN(n6132) );
  DFFRX1 \CACHE_reg[0][147]  ( .D(n4893), .CK(clk), .RN(n478), .Q(
        \CACHE[0][147] ), .QN(n6133) );
  DFFRX1 \CACHE_reg[0][146]  ( .D(n4894), .CK(clk), .RN(n479), .Q(
        \CACHE[0][146] ), .QN(n6134) );
  DFFRX1 \CACHE_reg[0][145]  ( .D(n4895), .CK(clk), .RN(n479), .Q(
        \CACHE[0][145] ), .QN(n6135) );
  DFFRX1 \CACHE_reg[0][144]  ( .D(n4896), .CK(clk), .RN(n480), .Q(
        \CACHE[0][144] ), .QN(n6136) );
  DFFRX1 \CACHE_reg[0][143]  ( .D(n4897), .CK(clk), .RN(n481), .Q(
        \CACHE[0][143] ), .QN(n6137) );
  DFFRX1 \CACHE_reg[0][142]  ( .D(n4898), .CK(clk), .RN(n481), .Q(
        \CACHE[0][142] ), .QN(n6138) );
  DFFRX1 \CACHE_reg[0][141]  ( .D(n4899), .CK(clk), .RN(n482), .Q(
        \CACHE[0][141] ), .QN(n6139) );
  DFFRX1 \CACHE_reg[0][140]  ( .D(n4900), .CK(clk), .RN(n483), .Q(
        \CACHE[0][140] ), .QN(n6140) );
  DFFRX1 \CACHE_reg[0][139]  ( .D(n4901), .CK(clk), .RN(n490), .Q(
        \CACHE[0][139] ), .QN(n6141) );
  DFFRX1 \CACHE_reg[0][138]  ( .D(n4902), .CK(clk), .RN(n483), .Q(
        \CACHE[0][138] ), .QN(n6142) );
  DFFRX1 \CACHE_reg[0][137]  ( .D(n4903), .CK(clk), .RN(n484), .Q(
        \CACHE[0][137] ), .QN(n6143) );
  DFFRX1 \CACHE_reg[0][136]  ( .D(n4904), .CK(clk), .RN(n485), .Q(
        \CACHE[0][136] ), .QN(n6144) );
  DFFRX1 \CACHE_reg[0][135]  ( .D(n4905), .CK(clk), .RN(n485), .Q(
        \CACHE[0][135] ), .QN(n6145) );
  DFFRX1 \CACHE_reg[0][134]  ( .D(n4906), .CK(clk), .RN(n486), .Q(
        \CACHE[0][134] ), .QN(n6146) );
  DFFRX1 \CACHE_reg[0][133]  ( .D(n4907), .CK(clk), .RN(n487), .Q(
        \CACHE[0][133] ), .QN(n6147) );
  DFFRX1 \CACHE_reg[0][132]  ( .D(n4908), .CK(clk), .RN(n474), .Q(
        \CACHE[0][132] ), .QN(n6148) );
  DFFRX1 \CACHE_reg[0][131]  ( .D(n4909), .CK(clk), .RN(n487), .Q(
        \CACHE[0][131] ), .QN(n6149) );
  DFFRX1 \CACHE_reg[0][130]  ( .D(n4910), .CK(clk), .RN(n488), .Q(
        \CACHE[0][130] ), .QN(n6150) );
  DFFRX1 \CACHE_reg[0][129]  ( .D(n4911), .CK(clk), .RN(n489), .Q(
        \CACHE[0][129] ), .QN(n6151) );
  DFFRX1 \CACHE_reg[0][128]  ( .D(n4912), .CK(clk), .RN(n489), .Q(
        \CACHE[0][128] ), .QN(n6152) );
  DFFRX1 \CACHE_reg[0][127]  ( .D(n4913), .CK(clk), .RN(n3056), .Q(
        \CACHE[0][127] ), .QN(n6153) );
  DFFRX1 \CACHE_reg[0][126]  ( .D(n4914), .CK(clk), .RN(n492), .Q(
        \CACHE[0][126] ), .QN(n6154) );
  DFFRX1 \CACHE_reg[0][125]  ( .D(n4915), .CK(clk), .RN(n534), .Q(
        \CACHE[0][125] ), .QN(n6155) );
  DFFRX1 \CACHE_reg[0][124]  ( .D(n4916), .CK(clk), .RN(n534), .Q(
        \CACHE[0][124] ), .QN(n6156) );
  DFFRX1 \CACHE_reg[0][123]  ( .D(n4917), .CK(clk), .RN(n535), .Q(
        \CACHE[0][123] ), .QN(n6157) );
  DFFRX1 \CACHE_reg[0][122]  ( .D(n4918), .CK(clk), .RN(n536), .Q(
        \CACHE[0][122] ), .QN(n6158) );
  DFFRX1 \CACHE_reg[0][121]  ( .D(n4919), .CK(clk), .RN(n536), .Q(
        \CACHE[0][121] ), .QN(n6159) );
  DFFRX1 \CACHE_reg[0][120]  ( .D(n4920), .CK(clk), .RN(n537), .Q(
        \CACHE[0][120] ), .QN(n6160) );
  DFFRX1 \CACHE_reg[0][119]  ( .D(n4921), .CK(clk), .RN(n538), .Q(
        \CACHE[0][119] ), .QN(n6161) );
  DFFRX1 \CACHE_reg[0][118]  ( .D(n4922), .CK(clk), .RN(n538), .Q(
        \CACHE[0][118] ), .QN(n6162) );
  DFFRX1 \CACHE_reg[0][117]  ( .D(n4923), .CK(clk), .RN(n539), .Q(
        \CACHE[0][117] ), .QN(n6163) );
  DFFRX1 \CACHE_reg[0][116]  ( .D(n4924), .CK(clk), .RN(n540), .Q(
        \CACHE[0][116] ), .QN(n6164) );
  DFFRX1 \CACHE_reg[0][115]  ( .D(n4925), .CK(clk), .RN(n540), .Q(
        \CACHE[0][115] ), .QN(n6165) );
  DFFRX1 \CACHE_reg[0][114]  ( .D(n4926), .CK(clk), .RN(n3020), .Q(
        \CACHE[0][114] ), .QN(n6166) );
  DFFRX1 \CACHE_reg[0][113]  ( .D(n4927), .CK(clk), .RN(n3022), .Q(
        \CACHE[0][113] ), .QN(n6167) );
  DFFRX1 \CACHE_reg[0][112]  ( .D(n4928), .CK(clk), .RN(n3022), .Q(
        \CACHE[0][112] ), .QN(n6168) );
  DFFRX1 \CACHE_reg[0][111]  ( .D(n4929), .CK(clk), .RN(n3023), .Q(
        \CACHE[0][111] ), .QN(n6169) );
  DFFRX1 \CACHE_reg[0][110]  ( .D(n4930), .CK(clk), .RN(n3024), .Q(
        \CACHE[0][110] ), .QN(n6170) );
  DFFRX1 \CACHE_reg[0][109]  ( .D(n4931), .CK(clk), .RN(n3024), .Q(
        \CACHE[0][109] ), .QN(n6171) );
  DFFRX1 \CACHE_reg[0][108]  ( .D(n4932), .CK(clk), .RN(n3025), .Q(
        \CACHE[0][108] ), .QN(n6172) );
  DFFRX1 \CACHE_reg[0][107]  ( .D(n4933), .CK(clk), .RN(n3026), .Q(
        \CACHE[0][107] ), .QN(n6173) );
  DFFRX1 \CACHE_reg[0][106]  ( .D(n4934), .CK(clk), .RN(n3026), .Q(
        \CACHE[0][106] ), .QN(n6174) );
  DFFRX1 \CACHE_reg[0][105]  ( .D(n4935), .CK(clk), .RN(n3027), .Q(
        \CACHE[0][105] ), .QN(n6175) );
  DFFRX1 \CACHE_reg[0][104]  ( .D(n4936), .CK(clk), .RN(n3028), .Q(
        \CACHE[0][104] ), .QN(n6176) );
  DFFRX1 \CACHE_reg[0][103]  ( .D(n4937), .CK(clk), .RN(n3028), .Q(
        \CACHE[0][103] ), .QN(n6177) );
  DFFRX1 \CACHE_reg[0][102]  ( .D(n4938), .CK(clk), .RN(n3029), .Q(
        \CACHE[0][102] ), .QN(n6178) );
  DFFRX1 \CACHE_reg[0][101]  ( .D(n4939), .CK(clk), .RN(n3030), .Q(
        \CACHE[0][101] ), .QN(n6179) );
  DFFRX1 \CACHE_reg[0][100]  ( .D(n4940), .CK(clk), .RN(n3030), .Q(
        \CACHE[0][100] ), .QN(n6180) );
  DFFRX1 \CACHE_reg[0][99]  ( .D(n4941), .CK(clk), .RN(n3031), .Q(
        \CACHE[0][99] ), .QN(n6181) );
  DFFRX1 \CACHE_reg[0][98]  ( .D(n4942), .CK(clk), .RN(n3032), .Q(
        \CACHE[0][98] ), .QN(n6182) );
  DFFRX1 \CACHE_reg[0][97]  ( .D(n4943), .CK(clk), .RN(n3032), .Q(
        \CACHE[0][97] ), .QN(n6183) );
  DFFRX1 \CACHE_reg[0][96]  ( .D(n4944), .CK(clk), .RN(n3033), .Q(
        \CACHE[0][96] ), .QN(n6184) );
  DFFRX1 \CACHE_reg[0][95]  ( .D(n4945), .CK(clk), .RN(n3034), .Q(
        \CACHE[0][95] ), .QN(n6185) );
  DFFRX1 \CACHE_reg[0][94]  ( .D(n4946), .CK(clk), .RN(n3034), .Q(
        \CACHE[0][94] ), .QN(n6186) );
  DFFRX1 \CACHE_reg[0][93]  ( .D(n4947), .CK(clk), .RN(n3035), .Q(
        \CACHE[0][93] ), .QN(n6187) );
  DFFRX1 \CACHE_reg[0][92]  ( .D(n4948), .CK(clk), .RN(n3036), .Q(
        \CACHE[0][92] ), .QN(n6188) );
  DFFRX1 \CACHE_reg[0][91]  ( .D(n4949), .CK(clk), .RN(n3036), .Q(
        \CACHE[0][91] ), .QN(n6189) );
  DFFRX1 \CACHE_reg[0][90]  ( .D(n4950), .CK(clk), .RN(n3037), .Q(
        \CACHE[0][90] ), .QN(n6190) );
  DFFRX1 \CACHE_reg[0][89]  ( .D(n4951), .CK(clk), .RN(n3038), .Q(
        \CACHE[0][89] ), .QN(n6191) );
  DFFRX1 \CACHE_reg[0][88]  ( .D(n4952), .CK(clk), .RN(n3038), .Q(
        \CACHE[0][88] ), .QN(n6192) );
  DFFRX1 \CACHE_reg[0][87]  ( .D(n4953), .CK(clk), .RN(n3039), .Q(
        \CACHE[0][87] ), .QN(n6193) );
  DFFRX1 \CACHE_reg[0][86]  ( .D(n4954), .CK(clk), .RN(n3040), .Q(
        \CACHE[0][86] ), .QN(n6194) );
  DFFRX1 \CACHE_reg[0][85]  ( .D(n4955), .CK(clk), .RN(n3040), .Q(
        \CACHE[0][85] ), .QN(n6195) );
  DFFRX1 \CACHE_reg[0][84]  ( .D(n4956), .CK(clk), .RN(n3041), .Q(
        \CACHE[0][84] ), .QN(n6196) );
  DFFRX1 \CACHE_reg[0][83]  ( .D(n4957), .CK(clk), .RN(n3042), .Q(
        \CACHE[0][83] ), .QN(n6197) );
  DFFRX1 \CACHE_reg[0][82]  ( .D(n4958), .CK(clk), .RN(n3042), .Q(
        \CACHE[0][82] ), .QN(n6198) );
  DFFRX1 \CACHE_reg[0][81]  ( .D(n4959), .CK(clk), .RN(n3043), .Q(
        \CACHE[0][81] ), .QN(n6199) );
  DFFRX1 \CACHE_reg[0][80]  ( .D(n4960), .CK(clk), .RN(n3044), .Q(
        \CACHE[0][80] ), .QN(n6200) );
  DFFRX1 \CACHE_reg[0][79]  ( .D(n4961), .CK(clk), .RN(n3044), .Q(
        \CACHE[0][79] ), .QN(n6201) );
  DFFRX1 \CACHE_reg[0][78]  ( .D(n4962), .CK(clk), .RN(n3045), .Q(
        \CACHE[0][78] ), .QN(n6202) );
  DFFRX1 \CACHE_reg[0][77]  ( .D(n4963), .CK(clk), .RN(n3046), .Q(
        \CACHE[0][77] ), .QN(n6203) );
  DFFRX1 \CACHE_reg[0][76]  ( .D(n4964), .CK(clk), .RN(n3046), .Q(
        \CACHE[0][76] ), .QN(n6204) );
  DFFRX1 \CACHE_reg[0][75]  ( .D(n4965), .CK(clk), .RN(n3047), .Q(
        \CACHE[0][75] ), .QN(n6205) );
  DFFRX1 \CACHE_reg[0][74]  ( .D(n4966), .CK(clk), .RN(n3048), .Q(
        \CACHE[0][74] ), .QN(n6206) );
  DFFRX1 \CACHE_reg[0][73]  ( .D(n4967), .CK(clk), .RN(n3048), .Q(
        \CACHE[0][73] ), .QN(n6207) );
  DFFRX1 \CACHE_reg[0][72]  ( .D(n4968), .CK(clk), .RN(n3049), .Q(
        \CACHE[0][72] ), .QN(n6208) );
  DFFRX1 \CACHE_reg[0][71]  ( .D(n4969), .CK(clk), .RN(n3050), .Q(
        \CACHE[0][71] ), .QN(n6209) );
  DFFRX1 \CACHE_reg[0][70]  ( .D(n4970), .CK(clk), .RN(n3050), .Q(
        \CACHE[0][70] ), .QN(n6210) );
  DFFRX1 \CACHE_reg[0][69]  ( .D(n4971), .CK(clk), .RN(n3051), .Q(
        \CACHE[0][69] ), .QN(n6211) );
  DFFRX1 \CACHE_reg[0][68]  ( .D(n4972), .CK(clk), .RN(n3052), .Q(
        \CACHE[0][68] ), .QN(n6212) );
  DFFRX1 \CACHE_reg[0][67]  ( .D(n4973), .CK(clk), .RN(n3052), .Q(
        \CACHE[0][67] ), .QN(n6213) );
  DFFRX1 \CACHE_reg[0][66]  ( .D(n4974), .CK(clk), .RN(n3053), .Q(
        \CACHE[0][66] ), .QN(n6214) );
  DFFRX1 \CACHE_reg[0][65]  ( .D(n4975), .CK(clk), .RN(n3054), .Q(
        \CACHE[0][65] ), .QN(n6215) );
  DFFRX1 \CACHE_reg[0][64]  ( .D(n4976), .CK(clk), .RN(n3054), .Q(
        \CACHE[0][64] ), .QN(n6216) );
  DFFRX1 \CACHE_reg[0][63]  ( .D(n4977), .CK(clk), .RN(n513), .Q(
        \CACHE[0][63] ), .QN(n6217) );
  DFFRX1 \CACHE_reg[0][62]  ( .D(n4978), .CK(clk), .RN(n513), .Q(
        \CACHE[0][62] ), .QN(n6218) );
  DFFRX1 \CACHE_reg[0][61]  ( .D(n4979), .CK(clk), .RN(n514), .Q(
        \CACHE[0][61] ), .QN(n6219) );
  DFFRX1 \CACHE_reg[0][60]  ( .D(n4980), .CK(clk), .RN(n515), .Q(
        \CACHE[0][60] ), .QN(n6220) );
  DFFRX1 \CACHE_reg[0][59]  ( .D(n4981), .CK(clk), .RN(n515), .Q(
        \CACHE[0][59] ), .QN(n6221) );
  DFFRX1 \CACHE_reg[0][58]  ( .D(n4982), .CK(clk), .RN(n516), .Q(
        \CACHE[0][58] ), .QN(n6222) );
  DFFRX1 \CACHE_reg[0][57]  ( .D(n4983), .CK(clk), .RN(n517), .Q(
        \CACHE[0][57] ), .QN(n6223) );
  DFFRX1 \CACHE_reg[0][56]  ( .D(n4984), .CK(clk), .RN(n517), .Q(
        \CACHE[0][56] ), .QN(n6224) );
  DFFRX1 \CACHE_reg[0][55]  ( .D(n4985), .CK(clk), .RN(n518), .Q(
        \CACHE[0][55] ), .QN(n6225) );
  DFFRX1 \CACHE_reg[0][54]  ( .D(n4986), .CK(clk), .RN(n519), .Q(
        \CACHE[0][54] ), .QN(n6226) );
  DFFRX1 \CACHE_reg[0][53]  ( .D(n4987), .CK(clk), .RN(n519), .Q(
        \CACHE[0][53] ), .QN(n6227) );
  DFFRX1 \CACHE_reg[0][52]  ( .D(n4988), .CK(clk), .RN(n520), .Q(
        \CACHE[0][52] ), .QN(n6228) );
  DFFRX1 \CACHE_reg[0][51]  ( .D(n4989), .CK(clk), .RN(n521), .Q(
        \CACHE[0][51] ), .QN(n6229) );
  DFFRX1 \CACHE_reg[0][50]  ( .D(n4990), .CK(clk), .RN(n521), .Q(
        \CACHE[0][50] ), .QN(n6230) );
  DFFRX1 \CACHE_reg[0][49]  ( .D(n4991), .CK(clk), .RN(n522), .Q(
        \CACHE[0][49] ), .QN(n6231) );
  DFFRX1 \CACHE_reg[0][48]  ( .D(n4992), .CK(clk), .RN(n523), .Q(
        \CACHE[0][48] ), .QN(n6232) );
  DFFRX1 \CACHE_reg[0][47]  ( .D(n4993), .CK(clk), .RN(n523), .Q(
        \CACHE[0][47] ), .QN(n6233) );
  DFFRX1 \CACHE_reg[0][46]  ( .D(n4994), .CK(clk), .RN(n524), .Q(
        \CACHE[0][46] ), .QN(n6234) );
  DFFRX1 \CACHE_reg[0][45]  ( .D(n4995), .CK(clk), .RN(n525), .Q(
        \CACHE[0][45] ), .QN(n6235) );
  DFFRX1 \CACHE_reg[0][44]  ( .D(n4996), .CK(clk), .RN(n525), .Q(
        \CACHE[0][44] ), .QN(n6236) );
  DFFRX1 \CACHE_reg[0][43]  ( .D(n4997), .CK(clk), .RN(n526), .Q(
        \CACHE[0][43] ), .QN(n6237) );
  DFFRX1 \CACHE_reg[0][42]  ( .D(n4998), .CK(clk), .RN(n527), .Q(
        \CACHE[0][42] ), .QN(n6238) );
  DFFRX1 \CACHE_reg[0][41]  ( .D(n4999), .CK(clk), .RN(n527), .Q(
        \CACHE[0][41] ), .QN(n6239) );
  DFFRX1 \CACHE_reg[0][40]  ( .D(n5000), .CK(clk), .RN(n528), .Q(
        \CACHE[0][40] ), .QN(n6240) );
  DFFRX1 \CACHE_reg[0][39]  ( .D(n5001), .CK(clk), .RN(n529), .Q(
        \CACHE[0][39] ), .QN(n6241) );
  DFFRX1 \CACHE_reg[0][38]  ( .D(n5002), .CK(clk), .RN(n529), .Q(
        \CACHE[0][38] ), .QN(n6242) );
  DFFRX1 \CACHE_reg[0][37]  ( .D(n5003), .CK(clk), .RN(n530), .Q(
        \CACHE[0][37] ), .QN(n6243) );
  DFFRX1 \CACHE_reg[0][36]  ( .D(n5004), .CK(clk), .RN(n531), .Q(
        \CACHE[0][36] ), .QN(n6244) );
  DFFRX1 \CACHE_reg[0][35]  ( .D(n5005), .CK(clk), .RN(n531), .Q(
        \CACHE[0][35] ), .QN(n6245) );
  DFFRX1 \CACHE_reg[0][34]  ( .D(n5006), .CK(clk), .RN(n532), .Q(
        \CACHE[0][34] ), .QN(n6246) );
  DFFRX1 \CACHE_reg[0][33]  ( .D(n5007), .CK(clk), .RN(n533), .Q(
        \CACHE[0][33] ), .QN(n6247) );
  DFFRX1 \CACHE_reg[0][32]  ( .D(n5008), .CK(clk), .RN(n533), .Q(
        \CACHE[0][32] ), .QN(n6248) );
  DFFRX1 \CACHE_reg[0][31]  ( .D(n5009), .CK(clk), .RN(n491), .Q(
        \CACHE[0][31] ), .QN(n6249) );
  DFFRX1 \CACHE_reg[0][30]  ( .D(n5010), .CK(clk), .RN(n3056), .Q(
        \CACHE[0][30] ), .QN(n6250) );
  DFFRX1 \CACHE_reg[0][29]  ( .D(n5011), .CK(clk), .RN(n493), .Q(
        \CACHE[0][29] ), .QN(n6251) );
  DFFRX1 \CACHE_reg[0][28]  ( .D(n5012), .CK(clk), .RN(n493), .Q(
        \CACHE[0][28] ), .QN(n6252) );
  DFFRX1 \CACHE_reg[0][27]  ( .D(n5013), .CK(clk), .RN(n494), .Q(
        \CACHE[0][27] ), .QN(n6253) );
  DFFRX1 \CACHE_reg[0][26]  ( .D(n5014), .CK(clk), .RN(n495), .Q(
        \CACHE[0][26] ), .QN(n6254) );
  DFFRX1 \CACHE_reg[0][25]  ( .D(n5015), .CK(clk), .RN(n495), .Q(
        \CACHE[0][25] ), .QN(n6255) );
  DFFRX1 \CACHE_reg[0][24]  ( .D(n5016), .CK(clk), .RN(n496), .Q(
        \CACHE[0][24] ), .QN(n6256) );
  DFFRX1 \CACHE_reg[0][23]  ( .D(n5017), .CK(clk), .RN(n497), .Q(
        \CACHE[0][23] ), .QN(n6257) );
  DFFRX1 \CACHE_reg[0][22]  ( .D(n5018), .CK(clk), .RN(n497), .Q(
        \CACHE[0][22] ), .QN(n6258) );
  DFFRX1 \CACHE_reg[0][21]  ( .D(n5019), .CK(clk), .RN(n498), .Q(
        \CACHE[0][21] ), .QN(n6259) );
  DFFRX1 \CACHE_reg[0][20]  ( .D(n5020), .CK(clk), .RN(n499), .Q(
        \CACHE[0][20] ), .QN(n6260) );
  DFFRX1 \CACHE_reg[0][19]  ( .D(n5021), .CK(clk), .RN(n499), .Q(
        \CACHE[0][19] ), .QN(n6261) );
  DFFRX1 \CACHE_reg[0][18]  ( .D(n5022), .CK(clk), .RN(n500), .Q(
        \CACHE[0][18] ), .QN(n6262) );
  DFFRX1 \CACHE_reg[0][17]  ( .D(n5023), .CK(clk), .RN(n501), .Q(
        \CACHE[0][17] ), .QN(n6263) );
  DFFRX1 \CACHE_reg[0][16]  ( .D(n5024), .CK(clk), .RN(n501), .Q(
        \CACHE[0][16] ), .QN(n6264) );
  DFFRX1 \CACHE_reg[0][15]  ( .D(n5025), .CK(clk), .RN(n502), .Q(
        \CACHE[0][15] ), .QN(n6265) );
  DFFRX1 \CACHE_reg[0][14]  ( .D(n5026), .CK(clk), .RN(n503), .Q(
        \CACHE[0][14] ), .QN(n6266) );
  DFFRX1 \CACHE_reg[0][13]  ( .D(n5027), .CK(clk), .RN(n503), .Q(
        \CACHE[0][13] ), .QN(n6267) );
  DFFRX1 \CACHE_reg[0][12]  ( .D(n5028), .CK(clk), .RN(n504), .Q(
        \CACHE[0][12] ), .QN(n6268) );
  DFFRX1 \CACHE_reg[0][11]  ( .D(n5029), .CK(clk), .RN(n505), .Q(
        \CACHE[0][11] ), .QN(n6269) );
  DFFRX1 \CACHE_reg[0][10]  ( .D(n5030), .CK(clk), .RN(n505), .Q(
        \CACHE[0][10] ), .QN(n6270) );
  DFFRX1 \CACHE_reg[0][9]  ( .D(n5031), .CK(clk), .RN(n506), .Q(\CACHE[0][9] ), 
        .QN(n6271) );
  DFFRX1 \CACHE_reg[0][8]  ( .D(n5032), .CK(clk), .RN(n507), .Q(\CACHE[0][8] ), 
        .QN(n6272) );
  DFFRX1 \CACHE_reg[0][7]  ( .D(n5033), .CK(clk), .RN(n507), .Q(\CACHE[0][7] ), 
        .QN(n6273) );
  DFFRX1 \CACHE_reg[0][6]  ( .D(n5034), .CK(clk), .RN(n508), .Q(\CACHE[0][6] ), 
        .QN(n6274) );
  DFFRX1 \CACHE_reg[0][5]  ( .D(n5035), .CK(clk), .RN(n509), .Q(\CACHE[0][5] ), 
        .QN(n6275) );
  DFFRX1 \CACHE_reg[0][4]  ( .D(n5036), .CK(clk), .RN(n509), .Q(\CACHE[0][4] ), 
        .QN(n6276) );
  DFFRX1 \CACHE_reg[0][3]  ( .D(n5037), .CK(clk), .RN(n510), .Q(\CACHE[0][3] ), 
        .QN(n6277) );
  DFFRX1 \CACHE_reg[0][2]  ( .D(n5038), .CK(clk), .RN(n511), .Q(\CACHE[0][2] ), 
        .QN(n6278) );
  DFFRX1 \CACHE_reg[0][1]  ( .D(n5039), .CK(clk), .RN(n511), .Q(\CACHE[0][1] ), 
        .QN(n6279) );
  DFFRX1 \CACHE_reg[0][0]  ( .D(n5040), .CK(clk), .RN(n512), .Q(\CACHE[0][0] ), 
        .QN(n6280) );
  DFFRX1 \CACHE_reg[6][154]  ( .D(n3956), .CK(clk), .RN(n491), .Q(
        \CACHE[6][154] ), .QN(n5196) );
  DFFRX1 \CACHE_reg[6][153]  ( .D(n3957), .CK(clk), .RN(n491), .Q(
        \CACHE[6][153] ), .QN(n5197) );
  DFFRX1 \CACHE_reg[6][152]  ( .D(n3958), .CK(clk), .RN(n474), .Q(
        \CACHE[6][152] ), .QN(n5198) );
  DFFRX1 \CACHE_reg[6][151]  ( .D(n3959), .CK(clk), .RN(n475), .Q(
        \CACHE[6][151] ), .QN(n5199) );
  DFFRX1 \CACHE_reg[6][150]  ( .D(n3960), .CK(clk), .RN(n476), .Q(
        \CACHE[6][150] ), .QN(n5200) );
  DFFRX1 \CACHE_reg[6][149]  ( .D(n3961), .CK(clk), .RN(n476), .Q(
        \CACHE[6][149] ), .QN(n5201) );
  DFFRX1 \CACHE_reg[6][148]  ( .D(n3962), .CK(clk), .RN(n477), .Q(
        \CACHE[6][148] ), .QN(n5202) );
  DFFRX1 \CACHE_reg[6][147]  ( .D(n3963), .CK(clk), .RN(n478), .Q(
        \CACHE[6][147] ), .QN(n5203) );
  DFFRX1 \CACHE_reg[6][146]  ( .D(n3964), .CK(clk), .RN(n478), .Q(
        \CACHE[6][146] ), .QN(n5204) );
  DFFRX1 \CACHE_reg[6][145]  ( .D(n3965), .CK(clk), .RN(n479), .Q(
        \CACHE[6][145] ), .QN(n5205) );
  DFFRX1 \CACHE_reg[6][144]  ( .D(n3966), .CK(clk), .RN(n480), .Q(
        \CACHE[6][144] ), .QN(n5206) );
  DFFRX1 \CACHE_reg[6][143]  ( .D(n3967), .CK(clk), .RN(n480), .Q(
        \CACHE[6][143] ), .QN(n5207) );
  DFFRX1 \CACHE_reg[6][142]  ( .D(n3968), .CK(clk), .RN(n481), .Q(
        \CACHE[6][142] ), .QN(n5208) );
  DFFRX1 \CACHE_reg[6][141]  ( .D(n3969), .CK(clk), .RN(n482), .Q(
        \CACHE[6][141] ), .QN(n5209) );
  DFFRX1 \CACHE_reg[6][140]  ( .D(n3970), .CK(clk), .RN(n482), .Q(
        \CACHE[6][140] ), .QN(n5210) );
  DFFRX1 \CACHE_reg[6][139]  ( .D(n3971), .CK(clk), .RN(n490), .Q(
        \CACHE[6][139] ), .QN(n5211) );
  DFFRX1 \CACHE_reg[6][138]  ( .D(n3972), .CK(clk), .RN(n483), .Q(
        \CACHE[6][138] ), .QN(n5212) );
  DFFRX1 \CACHE_reg[6][137]  ( .D(n3973), .CK(clk), .RN(n484), .Q(
        \CACHE[6][137] ), .QN(n5213) );
  DFFRX1 \CACHE_reg[6][136]  ( .D(n3974), .CK(clk), .RN(n484), .Q(
        \CACHE[6][136] ), .QN(n5214) );
  DFFRX1 \CACHE_reg[6][135]  ( .D(n3975), .CK(clk), .RN(n485), .Q(
        \CACHE[6][135] ), .QN(n5215) );
  DFFRX1 \CACHE_reg[6][134]  ( .D(n3976), .CK(clk), .RN(n486), .Q(
        \CACHE[6][134] ), .QN(n5216) );
  DFFRX1 \CACHE_reg[6][133]  ( .D(n3977), .CK(clk), .RN(n486), .Q(
        \CACHE[6][133] ), .QN(n5217) );
  DFFRX1 \CACHE_reg[6][132]  ( .D(n3978), .CK(clk), .RN(n474), .Q(
        \CACHE[6][132] ), .QN(n5218) );
  DFFRX1 \CACHE_reg[6][131]  ( .D(n3979), .CK(clk), .RN(n487), .Q(
        \CACHE[6][131] ), .QN(n5219) );
  DFFRX1 \CACHE_reg[6][130]  ( .D(n3980), .CK(clk), .RN(n488), .Q(
        \CACHE[6][130] ), .QN(n5220) );
  DFFRX1 \CACHE_reg[6][129]  ( .D(n3981), .CK(clk), .RN(n488), .Q(
        \CACHE[6][129] ), .QN(n5221) );
  DFFRX1 \CACHE_reg[6][128]  ( .D(n3982), .CK(clk), .RN(n489), .Q(
        \CACHE[6][128] ), .QN(n5222) );
  DFFRX1 \CACHE_reg[6][127]  ( .D(n3983), .CK(clk), .RN(n491), .Q(
        \CACHE[6][127] ), .QN(n5223) );
  DFFRX1 \CACHE_reg[6][126]  ( .D(n3984), .CK(clk), .RN(n492), .Q(
        \CACHE[6][126] ), .QN(n5224) );
  DFFRX1 \CACHE_reg[6][125]  ( .D(n3985), .CK(clk), .RN(n3056), .Q(
        \CACHE[6][125] ), .QN(n5225) );
  DFFRX1 \CACHE_reg[6][124]  ( .D(n3986), .CK(clk), .RN(n534), .Q(
        \CACHE[6][124] ), .QN(n5226) );
  DFFRX1 \CACHE_reg[6][123]  ( .D(n3987), .CK(clk), .RN(n535), .Q(
        \CACHE[6][123] ), .QN(n5227) );
  DFFRX1 \CACHE_reg[6][122]  ( .D(n3988), .CK(clk), .RN(n535), .Q(
        \CACHE[6][122] ), .QN(n5228) );
  DFFRX1 \CACHE_reg[6][121]  ( .D(n3989), .CK(clk), .RN(n536), .Q(
        \CACHE[6][121] ), .QN(n5229) );
  DFFRX1 \CACHE_reg[6][120]  ( .D(n3990), .CK(clk), .RN(n537), .Q(
        \CACHE[6][120] ), .QN(n5230) );
  DFFRX1 \CACHE_reg[6][119]  ( .D(n3991), .CK(clk), .RN(n537), .Q(
        \CACHE[6][119] ), .QN(n5231) );
  DFFRX1 \CACHE_reg[6][118]  ( .D(n3992), .CK(clk), .RN(n538), .Q(
        \CACHE[6][118] ), .QN(n5232) );
  DFFRX1 \CACHE_reg[6][117]  ( .D(n3993), .CK(clk), .RN(n539), .Q(
        \CACHE[6][117] ), .QN(n5233) );
  DFFRX1 \CACHE_reg[6][116]  ( .D(n3994), .CK(clk), .RN(n539), .Q(
        \CACHE[6][116] ), .QN(n5234) );
  DFFRX1 \CACHE_reg[6][115]  ( .D(n3995), .CK(clk), .RN(n540), .Q(
        \CACHE[6][115] ), .QN(n5235) );
  DFFRX1 \CACHE_reg[6][114]  ( .D(n3996), .CK(clk), .RN(n3020), .Q(
        \CACHE[6][114] ), .QN(n5236) );
  DFFRX1 \CACHE_reg[6][113]  ( .D(n3997), .CK(clk), .RN(n3020), .Q(
        \CACHE[6][113] ), .QN(n5237) );
  DFFRX1 \CACHE_reg[6][112]  ( .D(n3998), .CK(clk), .RN(n3022), .Q(
        \CACHE[6][112] ), .QN(n5238) );
  DFFRX1 \CACHE_reg[6][111]  ( .D(n3999), .CK(clk), .RN(n3023), .Q(
        \CACHE[6][111] ), .QN(n5239) );
  DFFRX1 \CACHE_reg[6][110]  ( .D(n4000), .CK(clk), .RN(n3023), .Q(
        \CACHE[6][110] ), .QN(n5240) );
  DFFRX1 \CACHE_reg[6][109]  ( .D(n4001), .CK(clk), .RN(n3024), .Q(
        \CACHE[6][109] ), .QN(n5241) );
  DFFRX1 \CACHE_reg[6][108]  ( .D(n4002), .CK(clk), .RN(n3025), .Q(
        \CACHE[6][108] ), .QN(n5242) );
  DFFRX1 \CACHE_reg[6][107]  ( .D(n4003), .CK(clk), .RN(n3025), .Q(
        \CACHE[6][107] ), .QN(n5243) );
  DFFRX1 \CACHE_reg[6][106]  ( .D(n4004), .CK(clk), .RN(n3026), .Q(
        \CACHE[6][106] ), .QN(n5244) );
  DFFRX1 \CACHE_reg[6][105]  ( .D(n4005), .CK(clk), .RN(n3027), .Q(
        \CACHE[6][105] ), .QN(n5245) );
  DFFRX1 \CACHE_reg[6][104]  ( .D(n4006), .CK(clk), .RN(n3027), .Q(
        \CACHE[6][104] ), .QN(n5246) );
  DFFRX1 \CACHE_reg[6][103]  ( .D(n4007), .CK(clk), .RN(n3028), .Q(
        \CACHE[6][103] ), .QN(n5247) );
  DFFRX1 \CACHE_reg[6][102]  ( .D(n4008), .CK(clk), .RN(n3029), .Q(
        \CACHE[6][102] ), .QN(n5248) );
  DFFRX1 \CACHE_reg[6][101]  ( .D(n4009), .CK(clk), .RN(n3029), .Q(
        \CACHE[6][101] ), .QN(n5249) );
  DFFRX1 \CACHE_reg[6][100]  ( .D(n4010), .CK(clk), .RN(n3030), .Q(
        \CACHE[6][100] ), .QN(n5250) );
  DFFRX1 \CACHE_reg[6][99]  ( .D(n4011), .CK(clk), .RN(n3031), .Q(
        \CACHE[6][99] ), .QN(n5251) );
  DFFRX1 \CACHE_reg[6][98]  ( .D(n4012), .CK(clk), .RN(n3031), .Q(
        \CACHE[6][98] ), .QN(n5252) );
  DFFRX1 \CACHE_reg[6][97]  ( .D(n4013), .CK(clk), .RN(n3032), .Q(
        \CACHE[6][97] ), .QN(n5253) );
  DFFRX1 \CACHE_reg[6][96]  ( .D(n4014), .CK(clk), .RN(n3033), .Q(
        \CACHE[6][96] ), .QN(n5254) );
  DFFRX1 \CACHE_reg[6][95]  ( .D(n4015), .CK(clk), .RN(n3033), .Q(
        \CACHE[6][95] ), .QN(n5255) );
  DFFRX1 \CACHE_reg[6][94]  ( .D(n4016), .CK(clk), .RN(n3034), .Q(
        \CACHE[6][94] ), .QN(n5256) );
  DFFRX1 \CACHE_reg[6][93]  ( .D(n4017), .CK(clk), .RN(n3035), .Q(
        \CACHE[6][93] ), .QN(n5257) );
  DFFRX1 \CACHE_reg[6][92]  ( .D(n4018), .CK(clk), .RN(n3035), .Q(
        \CACHE[6][92] ), .QN(n5258) );
  DFFRX1 \CACHE_reg[6][91]  ( .D(n4019), .CK(clk), .RN(n3036), .Q(
        \CACHE[6][91] ), .QN(n5259) );
  DFFRX1 \CACHE_reg[6][90]  ( .D(n4020), .CK(clk), .RN(n3037), .Q(
        \CACHE[6][90] ), .QN(n5260) );
  DFFRX1 \CACHE_reg[6][89]  ( .D(n4021), .CK(clk), .RN(n3037), .Q(
        \CACHE[6][89] ), .QN(n5261) );
  DFFRX1 \CACHE_reg[6][88]  ( .D(n4022), .CK(clk), .RN(n3038), .Q(
        \CACHE[6][88] ), .QN(n5262) );
  DFFRX1 \CACHE_reg[6][87]  ( .D(n4023), .CK(clk), .RN(n3039), .Q(
        \CACHE[6][87] ), .QN(n5263) );
  DFFRX1 \CACHE_reg[6][86]  ( .D(n4024), .CK(clk), .RN(n3039), .Q(
        \CACHE[6][86] ), .QN(n5264) );
  DFFRX1 \CACHE_reg[6][85]  ( .D(n4025), .CK(clk), .RN(n3040), .Q(
        \CACHE[6][85] ), .QN(n5265) );
  DFFRX1 \CACHE_reg[6][84]  ( .D(n4026), .CK(clk), .RN(n3041), .Q(
        \CACHE[6][84] ), .QN(n5266) );
  DFFRX1 \CACHE_reg[6][83]  ( .D(n4027), .CK(clk), .RN(n3041), .Q(
        \CACHE[6][83] ), .QN(n5267) );
  DFFRX1 \CACHE_reg[6][82]  ( .D(n4028), .CK(clk), .RN(n3042), .Q(
        \CACHE[6][82] ), .QN(n5268) );
  DFFRX1 \CACHE_reg[6][81]  ( .D(n4029), .CK(clk), .RN(n3043), .Q(
        \CACHE[6][81] ), .QN(n5269) );
  DFFRX1 \CACHE_reg[6][80]  ( .D(n4030), .CK(clk), .RN(n3043), .Q(
        \CACHE[6][80] ), .QN(n5270) );
  DFFRX1 \CACHE_reg[6][79]  ( .D(n4031), .CK(clk), .RN(n3044), .Q(
        \CACHE[6][79] ), .QN(n5271) );
  DFFRX1 \CACHE_reg[6][78]  ( .D(n4032), .CK(clk), .RN(n3045), .Q(
        \CACHE[6][78] ), .QN(n5272) );
  DFFRX1 \CACHE_reg[6][77]  ( .D(n4033), .CK(clk), .RN(n3045), .Q(
        \CACHE[6][77] ), .QN(n5273) );
  DFFRX1 \CACHE_reg[6][76]  ( .D(n4034), .CK(clk), .RN(n3046), .Q(
        \CACHE[6][76] ), .QN(n5274) );
  DFFRX1 \CACHE_reg[6][75]  ( .D(n4035), .CK(clk), .RN(n3047), .Q(
        \CACHE[6][75] ), .QN(n5275) );
  DFFRX1 \CACHE_reg[6][74]  ( .D(n4036), .CK(clk), .RN(n3047), .Q(
        \CACHE[6][74] ), .QN(n5276) );
  DFFRX1 \CACHE_reg[6][73]  ( .D(n4037), .CK(clk), .RN(n3048), .Q(
        \CACHE[6][73] ), .QN(n5277) );
  DFFRX1 \CACHE_reg[6][72]  ( .D(n4038), .CK(clk), .RN(n3049), .Q(
        \CACHE[6][72] ), .QN(n5278) );
  DFFRX1 \CACHE_reg[6][71]  ( .D(n4039), .CK(clk), .RN(n3049), .Q(
        \CACHE[6][71] ), .QN(n5279) );
  DFFRX1 \CACHE_reg[6][70]  ( .D(n4040), .CK(clk), .RN(n3050), .Q(
        \CACHE[6][70] ), .QN(n5280) );
  DFFRX1 \CACHE_reg[6][69]  ( .D(n4041), .CK(clk), .RN(n3051), .Q(
        \CACHE[6][69] ), .QN(n5281) );
  DFFRX1 \CACHE_reg[6][68]  ( .D(n4042), .CK(clk), .RN(n3051), .Q(
        \CACHE[6][68] ), .QN(n5282) );
  DFFRX1 \CACHE_reg[6][67]  ( .D(n4043), .CK(clk), .RN(n3052), .Q(
        \CACHE[6][67] ), .QN(n5283) );
  DFFRX1 \CACHE_reg[6][66]  ( .D(n4044), .CK(clk), .RN(n3053), .Q(
        \CACHE[6][66] ), .QN(n5284) );
  DFFRX1 \CACHE_reg[6][65]  ( .D(n4045), .CK(clk), .RN(n3053), .Q(
        \CACHE[6][65] ), .QN(n5285) );
  DFFRX1 \CACHE_reg[6][64]  ( .D(n4046), .CK(clk), .RN(n3054), .Q(
        \CACHE[6][64] ), .QN(n5286) );
  DFFRX1 \CACHE_reg[6][63]  ( .D(n4047), .CK(clk), .RN(n512), .Q(
        \CACHE[6][63] ), .QN(n5287) );
  DFFRX1 \CACHE_reg[6][62]  ( .D(n4048), .CK(clk), .RN(n513), .Q(
        \CACHE[6][62] ), .QN(n5288) );
  DFFRX1 \CACHE_reg[6][61]  ( .D(n4049), .CK(clk), .RN(n514), .Q(
        \CACHE[6][61] ), .QN(n5289) );
  DFFRX1 \CACHE_reg[6][60]  ( .D(n4050), .CK(clk), .RN(n514), .Q(
        \CACHE[6][60] ), .QN(n5290) );
  DFFRX1 \CACHE_reg[6][59]  ( .D(n4051), .CK(clk), .RN(n515), .Q(
        \CACHE[6][59] ), .QN(n5291) );
  DFFRX1 \CACHE_reg[6][58]  ( .D(n4052), .CK(clk), .RN(n516), .Q(
        \CACHE[6][58] ), .QN(n5292) );
  DFFRX1 \CACHE_reg[6][57]  ( .D(n4053), .CK(clk), .RN(n516), .Q(
        \CACHE[6][57] ), .QN(n5293) );
  DFFRX1 \CACHE_reg[6][56]  ( .D(n4054), .CK(clk), .RN(n517), .Q(
        \CACHE[6][56] ), .QN(n5294) );
  DFFRX1 \CACHE_reg[6][55]  ( .D(n4055), .CK(clk), .RN(n518), .Q(
        \CACHE[6][55] ), .QN(n5295) );
  DFFRX1 \CACHE_reg[6][54]  ( .D(n4056), .CK(clk), .RN(n518), .Q(
        \CACHE[6][54] ), .QN(n5296) );
  DFFRX1 \CACHE_reg[6][53]  ( .D(n4057), .CK(clk), .RN(n519), .Q(
        \CACHE[6][53] ), .QN(n5297) );
  DFFRX1 \CACHE_reg[6][52]  ( .D(n4058), .CK(clk), .RN(n520), .Q(
        \CACHE[6][52] ), .QN(n5298) );
  DFFRX1 \CACHE_reg[6][51]  ( .D(n4059), .CK(clk), .RN(n520), .Q(
        \CACHE[6][51] ), .QN(n5299) );
  DFFRX1 \CACHE_reg[6][50]  ( .D(n4060), .CK(clk), .RN(n521), .Q(
        \CACHE[6][50] ), .QN(n5300) );
  DFFRX1 \CACHE_reg[6][49]  ( .D(n4061), .CK(clk), .RN(n522), .Q(
        \CACHE[6][49] ), .QN(n5301) );
  DFFRX1 \CACHE_reg[6][48]  ( .D(n4062), .CK(clk), .RN(n522), .Q(
        \CACHE[6][48] ), .QN(n5302) );
  DFFRX1 \CACHE_reg[6][47]  ( .D(n4063), .CK(clk), .RN(n523), .Q(
        \CACHE[6][47] ), .QN(n5303) );
  DFFRX1 \CACHE_reg[6][46]  ( .D(n4064), .CK(clk), .RN(n524), .Q(
        \CACHE[6][46] ), .QN(n5304) );
  DFFRX1 \CACHE_reg[6][45]  ( .D(n4065), .CK(clk), .RN(n524), .Q(
        \CACHE[6][45] ), .QN(n5305) );
  DFFRX1 \CACHE_reg[6][44]  ( .D(n4066), .CK(clk), .RN(n525), .Q(
        \CACHE[6][44] ), .QN(n5306) );
  DFFRX1 \CACHE_reg[6][43]  ( .D(n4067), .CK(clk), .RN(n526), .Q(
        \CACHE[6][43] ), .QN(n5307) );
  DFFRX1 \CACHE_reg[6][42]  ( .D(n4068), .CK(clk), .RN(n526), .Q(
        \CACHE[6][42] ), .QN(n5308) );
  DFFRX1 \CACHE_reg[6][41]  ( .D(n4069), .CK(clk), .RN(n527), .Q(
        \CACHE[6][41] ), .QN(n5309) );
  DFFRX1 \CACHE_reg[6][40]  ( .D(n4070), .CK(clk), .RN(n528), .Q(
        \CACHE[6][40] ), .QN(n5310) );
  DFFRX1 \CACHE_reg[6][39]  ( .D(n4071), .CK(clk), .RN(n528), .Q(
        \CACHE[6][39] ), .QN(n5311) );
  DFFRX1 \CACHE_reg[6][38]  ( .D(n4072), .CK(clk), .RN(n529), .Q(
        \CACHE[6][38] ), .QN(n5312) );
  DFFRX1 \CACHE_reg[6][37]  ( .D(n4073), .CK(clk), .RN(n530), .Q(
        \CACHE[6][37] ), .QN(n5313) );
  DFFRX1 \CACHE_reg[6][36]  ( .D(n4074), .CK(clk), .RN(n530), .Q(
        \CACHE[6][36] ), .QN(n5314) );
  DFFRX1 \CACHE_reg[6][35]  ( .D(n4075), .CK(clk), .RN(n531), .Q(
        \CACHE[6][35] ), .QN(n5315) );
  DFFRX1 \CACHE_reg[6][34]  ( .D(n4076), .CK(clk), .RN(n532), .Q(
        \CACHE[6][34] ), .QN(n5316) );
  DFFRX1 \CACHE_reg[6][33]  ( .D(n4077), .CK(clk), .RN(n532), .Q(
        \CACHE[6][33] ), .QN(n5317) );
  DFFRX1 \CACHE_reg[6][32]  ( .D(n4078), .CK(clk), .RN(n533), .Q(
        \CACHE[6][32] ), .QN(n5318) );
  DFFRX1 \CACHE_reg[6][31]  ( .D(n4079), .CK(clk), .RN(n490), .Q(
        \CACHE[6][31] ), .QN(n5319) );
  DFFRX1 \CACHE_reg[6][30]  ( .D(n4080), .CK(clk), .RN(n3056), .Q(
        \CACHE[6][30] ), .QN(n5320) );
  DFFRX1 \CACHE_reg[6][29]  ( .D(n4081), .CK(clk), .RN(n492), .Q(
        \CACHE[6][29] ), .QN(n5321) );
  DFFRX1 \CACHE_reg[6][28]  ( .D(n4082), .CK(clk), .RN(n493), .Q(
        \CACHE[6][28] ), .QN(n5322) );
  DFFRX1 \CACHE_reg[6][27]  ( .D(n4083), .CK(clk), .RN(n494), .Q(
        \CACHE[6][27] ), .QN(n5323) );
  DFFRX1 \CACHE_reg[6][26]  ( .D(n4084), .CK(clk), .RN(n494), .Q(
        \CACHE[6][26] ), .QN(n5324) );
  DFFRX1 \CACHE_reg[6][25]  ( .D(n4085), .CK(clk), .RN(n495), .Q(
        \CACHE[6][25] ), .QN(n5325) );
  DFFRX1 \CACHE_reg[6][24]  ( .D(n4086), .CK(clk), .RN(n496), .Q(
        \CACHE[6][24] ), .QN(n5326) );
  DFFRX1 \CACHE_reg[6][23]  ( .D(n4087), .CK(clk), .RN(n496), .Q(
        \CACHE[6][23] ), .QN(n5327) );
  DFFRX1 \CACHE_reg[6][22]  ( .D(n4088), .CK(clk), .RN(n497), .Q(
        \CACHE[6][22] ), .QN(n5328) );
  DFFRX1 \CACHE_reg[6][21]  ( .D(n4089), .CK(clk), .RN(n498), .Q(
        \CACHE[6][21] ), .QN(n5329) );
  DFFRX1 \CACHE_reg[6][20]  ( .D(n4090), .CK(clk), .RN(n498), .Q(
        \CACHE[6][20] ), .QN(n5330) );
  DFFRX1 \CACHE_reg[6][19]  ( .D(n4091), .CK(clk), .RN(n499), .Q(
        \CACHE[6][19] ), .QN(n5331) );
  DFFRX1 \CACHE_reg[6][18]  ( .D(n4092), .CK(clk), .RN(n500), .Q(
        \CACHE[6][18] ), .QN(n5332) );
  DFFRX1 \CACHE_reg[6][17]  ( .D(n4093), .CK(clk), .RN(n500), .Q(
        \CACHE[6][17] ), .QN(n5333) );
  DFFRX1 \CACHE_reg[6][16]  ( .D(n4094), .CK(clk), .RN(n501), .Q(
        \CACHE[6][16] ), .QN(n5334) );
  DFFRX1 \CACHE_reg[6][15]  ( .D(n4095), .CK(clk), .RN(n502), .Q(
        \CACHE[6][15] ), .QN(n5335) );
  DFFRX1 \CACHE_reg[6][14]  ( .D(n4096), .CK(clk), .RN(n502), .Q(
        \CACHE[6][14] ), .QN(n5336) );
  DFFRX1 \CACHE_reg[6][13]  ( .D(n4097), .CK(clk), .RN(n503), .Q(
        \CACHE[6][13] ), .QN(n5337) );
  DFFRX1 \CACHE_reg[6][12]  ( .D(n4098), .CK(clk), .RN(n504), .Q(
        \CACHE[6][12] ), .QN(n5338) );
  DFFRX1 \CACHE_reg[6][11]  ( .D(n4099), .CK(clk), .RN(n504), .Q(
        \CACHE[6][11] ), .QN(n5339) );
  DFFRX1 \CACHE_reg[6][10]  ( .D(n4100), .CK(clk), .RN(n505), .Q(
        \CACHE[6][10] ), .QN(n5340) );
  DFFRX1 \CACHE_reg[6][9]  ( .D(n4101), .CK(clk), .RN(n506), .Q(\CACHE[6][9] ), 
        .QN(n5341) );
  DFFRX1 \CACHE_reg[6][8]  ( .D(n4102), .CK(clk), .RN(n506), .Q(\CACHE[6][8] ), 
        .QN(n5342) );
  DFFRX1 \CACHE_reg[6][7]  ( .D(n4103), .CK(clk), .RN(n507), .Q(\CACHE[6][7] ), 
        .QN(n5343) );
  DFFRX1 \CACHE_reg[6][6]  ( .D(n4104), .CK(clk), .RN(n508), .Q(\CACHE[6][6] ), 
        .QN(n5344) );
  DFFRX1 \CACHE_reg[6][5]  ( .D(n4105), .CK(clk), .RN(n508), .Q(\CACHE[6][5] ), 
        .QN(n5345) );
  DFFRX1 \CACHE_reg[6][4]  ( .D(n4106), .CK(clk), .RN(n509), .Q(\CACHE[6][4] ), 
        .QN(n5346) );
  DFFRX1 \CACHE_reg[6][3]  ( .D(n4107), .CK(clk), .RN(n510), .Q(\CACHE[6][3] ), 
        .QN(n5347) );
  DFFRX1 \CACHE_reg[6][2]  ( .D(n4108), .CK(clk), .RN(n510), .Q(\CACHE[6][2] ), 
        .QN(n5348) );
  DFFRX1 \CACHE_reg[6][1]  ( .D(n4109), .CK(clk), .RN(n511), .Q(\CACHE[6][1] ), 
        .QN(n5349) );
  DFFRX1 \CACHE_reg[6][0]  ( .D(n4110), .CK(clk), .RN(n512), .Q(\CACHE[6][0] ), 
        .QN(n5350) );
  DFFRX1 \CACHE_reg[2][154]  ( .D(n4576), .CK(clk), .RN(n3056), .Q(
        \CACHE[2][154] ), .QN(n5816) );
  DFFRX1 \CACHE_reg[2][153]  ( .D(n4577), .CK(clk), .RN(n3056), .Q(
        \CACHE[2][153] ), .QN(n5817) );
  DFFRX1 \CACHE_reg[2][152]  ( .D(n4578), .CK(clk), .RN(n475), .Q(
        \CACHE[2][152] ), .QN(n5818) );
  DFFRX1 \CACHE_reg[2][151]  ( .D(n4579), .CK(clk), .RN(n475), .Q(
        \CACHE[2][151] ), .QN(n5819) );
  DFFRX1 \CACHE_reg[2][150]  ( .D(n4580), .CK(clk), .RN(n476), .Q(
        \CACHE[2][150] ), .QN(n5820) );
  DFFRX1 \CACHE_reg[2][149]  ( .D(n4581), .CK(clk), .RN(n477), .Q(
        \CACHE[2][149] ), .QN(n5821) );
  DFFRX1 \CACHE_reg[2][148]  ( .D(n4582), .CK(clk), .RN(n477), .Q(
        \CACHE[2][148] ), .QN(n5822) );
  DFFRX1 \CACHE_reg[2][147]  ( .D(n4583), .CK(clk), .RN(n478), .Q(
        \CACHE[2][147] ), .QN(n5823) );
  DFFRX1 \CACHE_reg[2][146]  ( .D(n4584), .CK(clk), .RN(n479), .Q(
        \CACHE[2][146] ), .QN(n5824) );
  DFFRX1 \CACHE_reg[2][145]  ( .D(n4585), .CK(clk), .RN(n479), .Q(
        \CACHE[2][145] ), .QN(n5825) );
  DFFRX1 \CACHE_reg[2][144]  ( .D(n4586), .CK(clk), .RN(n480), .Q(
        \CACHE[2][144] ), .QN(n5826) );
  DFFRX1 \CACHE_reg[2][143]  ( .D(n4587), .CK(clk), .RN(n481), .Q(
        \CACHE[2][143] ), .QN(n5827) );
  DFFRX1 \CACHE_reg[2][142]  ( .D(n4588), .CK(clk), .RN(n481), .Q(
        \CACHE[2][142] ), .QN(n5828) );
  DFFRX1 \CACHE_reg[2][141]  ( .D(n4589), .CK(clk), .RN(n482), .Q(
        \CACHE[2][141] ), .QN(n5829) );
  DFFRX1 \CACHE_reg[2][140]  ( .D(n4590), .CK(clk), .RN(n483), .Q(
        \CACHE[2][140] ), .QN(n5830) );
  DFFRX1 \CACHE_reg[2][139]  ( .D(n4591), .CK(clk), .RN(n490), .Q(
        \CACHE[2][139] ), .QN(n5831) );
  DFFRX1 \CACHE_reg[2][138]  ( .D(n4592), .CK(clk), .RN(n483), .Q(
        \CACHE[2][138] ), .QN(n5832) );
  DFFRX1 \CACHE_reg[2][137]  ( .D(n4593), .CK(clk), .RN(n484), .Q(
        \CACHE[2][137] ), .QN(n5833) );
  DFFRX1 \CACHE_reg[2][136]  ( .D(n4594), .CK(clk), .RN(n485), .Q(
        \CACHE[2][136] ), .QN(n5834) );
  DFFRX1 \CACHE_reg[2][135]  ( .D(n4595), .CK(clk), .RN(n485), .Q(
        \CACHE[2][135] ), .QN(n5835) );
  DFFRX1 \CACHE_reg[2][134]  ( .D(n4596), .CK(clk), .RN(n486), .Q(
        \CACHE[2][134] ), .QN(n5836) );
  DFFRX1 \CACHE_reg[2][133]  ( .D(n4597), .CK(clk), .RN(n487), .Q(
        \CACHE[2][133] ), .QN(n5837) );
  DFFRX1 \CACHE_reg[2][132]  ( .D(n4598), .CK(clk), .RN(n474), .Q(
        \CACHE[2][132] ), .QN(n5838) );
  DFFRX1 \CACHE_reg[2][131]  ( .D(n4599), .CK(clk), .RN(n487), .Q(
        \CACHE[2][131] ), .QN(n5839) );
  DFFRX1 \CACHE_reg[2][130]  ( .D(n4600), .CK(clk), .RN(n488), .Q(
        \CACHE[2][130] ), .QN(n5840) );
  DFFRX1 \CACHE_reg[2][129]  ( .D(n4601), .CK(clk), .RN(n489), .Q(
        \CACHE[2][129] ), .QN(n5841) );
  DFFRX1 \CACHE_reg[2][128]  ( .D(n4602), .CK(clk), .RN(n489), .Q(
        \CACHE[2][128] ), .QN(n5842) );
  DFFRX1 \CACHE_reg[2][127]  ( .D(n4603), .CK(clk), .RN(n3056), .Q(
        \CACHE[2][127] ), .QN(n5843) );
  DFFRX1 \CACHE_reg[2][126]  ( .D(n4604), .CK(clk), .RN(n491), .Q(
        \CACHE[2][126] ), .QN(n5844) );
  DFFRX1 \CACHE_reg[2][125]  ( .D(n4605), .CK(clk), .RN(n534), .Q(
        \CACHE[2][125] ), .QN(n5845) );
  DFFRX1 \CACHE_reg[2][124]  ( .D(n4606), .CK(clk), .RN(n534), .Q(
        \CACHE[2][124] ), .QN(n5846) );
  DFFRX1 \CACHE_reg[2][123]  ( .D(n4607), .CK(clk), .RN(n535), .Q(
        \CACHE[2][123] ), .QN(n5847) );
  DFFRX1 \CACHE_reg[2][122]  ( .D(n4608), .CK(clk), .RN(n536), .Q(
        \CACHE[2][122] ), .QN(n5848) );
  DFFRX1 \CACHE_reg[2][121]  ( .D(n4609), .CK(clk), .RN(n536), .Q(
        \CACHE[2][121] ), .QN(n5849) );
  DFFRX1 \CACHE_reg[2][120]  ( .D(n4610), .CK(clk), .RN(n537), .Q(
        \CACHE[2][120] ), .QN(n5850) );
  DFFRX1 \CACHE_reg[2][119]  ( .D(n4611), .CK(clk), .RN(n538), .Q(
        \CACHE[2][119] ), .QN(n5851) );
  DFFRX1 \CACHE_reg[2][118]  ( .D(n4612), .CK(clk), .RN(n538), .Q(
        \CACHE[2][118] ), .QN(n5852) );
  DFFRX1 \CACHE_reg[2][117]  ( .D(n4613), .CK(clk), .RN(n539), .Q(
        \CACHE[2][117] ), .QN(n5853) );
  DFFRX1 \CACHE_reg[2][116]  ( .D(n4614), .CK(clk), .RN(n540), .Q(
        \CACHE[2][116] ), .QN(n5854) );
  DFFRX1 \CACHE_reg[2][115]  ( .D(n4615), .CK(clk), .RN(n540), .Q(
        \CACHE[2][115] ), .QN(n5855) );
  DFFRX1 \CACHE_reg[2][114]  ( .D(n4616), .CK(clk), .RN(n3020), .Q(
        \CACHE[2][114] ), .QN(n5856) );
  DFFRX1 \CACHE_reg[2][113]  ( .D(n4617), .CK(clk), .RN(n3022), .Q(
        \CACHE[2][113] ), .QN(n5857) );
  DFFRX1 \CACHE_reg[2][112]  ( .D(n4618), .CK(clk), .RN(n3022), .Q(
        \CACHE[2][112] ), .QN(n5858) );
  DFFRX1 \CACHE_reg[2][111]  ( .D(n4619), .CK(clk), .RN(n3023), .Q(
        \CACHE[2][111] ), .QN(n5859) );
  DFFRX1 \CACHE_reg[2][110]  ( .D(n4620), .CK(clk), .RN(n3024), .Q(
        \CACHE[2][110] ), .QN(n5860) );
  DFFRX1 \CACHE_reg[2][109]  ( .D(n4621), .CK(clk), .RN(n3024), .Q(
        \CACHE[2][109] ), .QN(n5861) );
  DFFRX1 \CACHE_reg[2][108]  ( .D(n4622), .CK(clk), .RN(n3025), .Q(
        \CACHE[2][108] ), .QN(n5862) );
  DFFRX1 \CACHE_reg[2][107]  ( .D(n4623), .CK(clk), .RN(n3026), .Q(
        \CACHE[2][107] ), .QN(n5863) );
  DFFRX1 \CACHE_reg[2][106]  ( .D(n4624), .CK(clk), .RN(n3026), .Q(
        \CACHE[2][106] ), .QN(n5864) );
  DFFRX1 \CACHE_reg[2][105]  ( .D(n4625), .CK(clk), .RN(n3027), .Q(
        \CACHE[2][105] ), .QN(n5865) );
  DFFRX1 \CACHE_reg[2][104]  ( .D(n4626), .CK(clk), .RN(n3028), .Q(
        \CACHE[2][104] ), .QN(n5866) );
  DFFRX1 \CACHE_reg[2][103]  ( .D(n4627), .CK(clk), .RN(n3028), .Q(
        \CACHE[2][103] ), .QN(n5867) );
  DFFRX1 \CACHE_reg[2][102]  ( .D(n4628), .CK(clk), .RN(n3029), .Q(
        \CACHE[2][102] ), .QN(n5868) );
  DFFRX1 \CACHE_reg[2][101]  ( .D(n4629), .CK(clk), .RN(n3030), .Q(
        \CACHE[2][101] ), .QN(n5869) );
  DFFRX1 \CACHE_reg[2][100]  ( .D(n4630), .CK(clk), .RN(n3030), .Q(
        \CACHE[2][100] ), .QN(n5870) );
  DFFRX1 \CACHE_reg[2][99]  ( .D(n4631), .CK(clk), .RN(n3031), .Q(
        \CACHE[2][99] ), .QN(n5871) );
  DFFRX1 \CACHE_reg[2][98]  ( .D(n4632), .CK(clk), .RN(n3032), .Q(
        \CACHE[2][98] ), .QN(n5872) );
  DFFRX1 \CACHE_reg[2][97]  ( .D(n4633), .CK(clk), .RN(n3032), .Q(
        \CACHE[2][97] ), .QN(n5873) );
  DFFRX1 \CACHE_reg[2][96]  ( .D(n4634), .CK(clk), .RN(n3033), .Q(
        \CACHE[2][96] ), .QN(n5874) );
  DFFRX1 \CACHE_reg[2][95]  ( .D(n4635), .CK(clk), .RN(n3034), .Q(
        \CACHE[2][95] ), .QN(n5875) );
  DFFRX1 \CACHE_reg[2][94]  ( .D(n4636), .CK(clk), .RN(n3034), .Q(
        \CACHE[2][94] ), .QN(n5876) );
  DFFRX1 \CACHE_reg[2][93]  ( .D(n4637), .CK(clk), .RN(n3035), .Q(
        \CACHE[2][93] ), .QN(n5877) );
  DFFRX1 \CACHE_reg[2][92]  ( .D(n4638), .CK(clk), .RN(n3036), .Q(
        \CACHE[2][92] ), .QN(n5878) );
  DFFRX1 \CACHE_reg[2][91]  ( .D(n4639), .CK(clk), .RN(n3036), .Q(
        \CACHE[2][91] ), .QN(n5879) );
  DFFRX1 \CACHE_reg[2][90]  ( .D(n4640), .CK(clk), .RN(n3037), .Q(
        \CACHE[2][90] ), .QN(n5880) );
  DFFRX1 \CACHE_reg[2][89]  ( .D(n4641), .CK(clk), .RN(n3038), .Q(
        \CACHE[2][89] ), .QN(n5881) );
  DFFRX1 \CACHE_reg[2][88]  ( .D(n4642), .CK(clk), .RN(n3038), .Q(
        \CACHE[2][88] ), .QN(n5882) );
  DFFRX1 \CACHE_reg[2][87]  ( .D(n4643), .CK(clk), .RN(n3039), .Q(
        \CACHE[2][87] ), .QN(n5883) );
  DFFRX1 \CACHE_reg[2][86]  ( .D(n4644), .CK(clk), .RN(n3040), .Q(
        \CACHE[2][86] ), .QN(n5884) );
  DFFRX1 \CACHE_reg[2][85]  ( .D(n4645), .CK(clk), .RN(n3040), .Q(
        \CACHE[2][85] ), .QN(n5885) );
  DFFRX1 \CACHE_reg[2][84]  ( .D(n4646), .CK(clk), .RN(n3041), .Q(
        \CACHE[2][84] ), .QN(n5886) );
  DFFRX1 \CACHE_reg[2][83]  ( .D(n4647), .CK(clk), .RN(n3042), .Q(
        \CACHE[2][83] ), .QN(n5887) );
  DFFRX1 \CACHE_reg[2][82]  ( .D(n4648), .CK(clk), .RN(n3042), .Q(
        \CACHE[2][82] ), .QN(n5888) );
  DFFRX1 \CACHE_reg[2][81]  ( .D(n4649), .CK(clk), .RN(n3043), .Q(
        \CACHE[2][81] ), .QN(n5889) );
  DFFRX1 \CACHE_reg[2][80]  ( .D(n4650), .CK(clk), .RN(n3044), .Q(
        \CACHE[2][80] ), .QN(n5890) );
  DFFRX1 \CACHE_reg[2][79]  ( .D(n4651), .CK(clk), .RN(n3044), .Q(
        \CACHE[2][79] ), .QN(n5891) );
  DFFRX1 \CACHE_reg[2][78]  ( .D(n4652), .CK(clk), .RN(n3045), .Q(
        \CACHE[2][78] ), .QN(n5892) );
  DFFRX1 \CACHE_reg[2][77]  ( .D(n4653), .CK(clk), .RN(n3046), .Q(
        \CACHE[2][77] ), .QN(n5893) );
  DFFRX1 \CACHE_reg[2][76]  ( .D(n4654), .CK(clk), .RN(n3046), .Q(
        \CACHE[2][76] ), .QN(n5894) );
  DFFRX1 \CACHE_reg[2][75]  ( .D(n4655), .CK(clk), .RN(n3047), .Q(
        \CACHE[2][75] ), .QN(n5895) );
  DFFRX1 \CACHE_reg[2][74]  ( .D(n4656), .CK(clk), .RN(n3048), .Q(
        \CACHE[2][74] ), .QN(n5896) );
  DFFRX1 \CACHE_reg[2][73]  ( .D(n4657), .CK(clk), .RN(n3048), .Q(
        \CACHE[2][73] ), .QN(n5897) );
  DFFRX1 \CACHE_reg[2][72]  ( .D(n4658), .CK(clk), .RN(n3049), .Q(
        \CACHE[2][72] ), .QN(n5898) );
  DFFRX1 \CACHE_reg[2][71]  ( .D(n4659), .CK(clk), .RN(n3050), .Q(
        \CACHE[2][71] ), .QN(n5899) );
  DFFRX1 \CACHE_reg[2][70]  ( .D(n4660), .CK(clk), .RN(n3050), .Q(
        \CACHE[2][70] ), .QN(n5900) );
  DFFRX1 \CACHE_reg[2][69]  ( .D(n4661), .CK(clk), .RN(n3051), .Q(
        \CACHE[2][69] ), .QN(n5901) );
  DFFRX1 \CACHE_reg[2][68]  ( .D(n4662), .CK(clk), .RN(n3052), .Q(
        \CACHE[2][68] ), .QN(n5902) );
  DFFRX1 \CACHE_reg[2][67]  ( .D(n4663), .CK(clk), .RN(n3052), .Q(
        \CACHE[2][67] ), .QN(n5903) );
  DFFRX1 \CACHE_reg[2][66]  ( .D(n4664), .CK(clk), .RN(n3053), .Q(
        \CACHE[2][66] ), .QN(n5904) );
  DFFRX1 \CACHE_reg[2][65]  ( .D(n4665), .CK(clk), .RN(n3054), .Q(
        \CACHE[2][65] ), .QN(n5905) );
  DFFRX1 \CACHE_reg[2][64]  ( .D(n4666), .CK(clk), .RN(n3054), .Q(
        \CACHE[2][64] ), .QN(n5906) );
  DFFRX1 \CACHE_reg[2][63]  ( .D(n4667), .CK(clk), .RN(n513), .Q(
        \CACHE[2][63] ), .QN(n5907) );
  DFFRX1 \CACHE_reg[2][62]  ( .D(n4668), .CK(clk), .RN(n513), .Q(
        \CACHE[2][62] ), .QN(n5908) );
  DFFRX1 \CACHE_reg[2][61]  ( .D(n4669), .CK(clk), .RN(n514), .Q(
        \CACHE[2][61] ), .QN(n5909) );
  DFFRX1 \CACHE_reg[2][60]  ( .D(n4670), .CK(clk), .RN(n515), .Q(
        \CACHE[2][60] ), .QN(n5910) );
  DFFRX1 \CACHE_reg[2][59]  ( .D(n4671), .CK(clk), .RN(n515), .Q(
        \CACHE[2][59] ), .QN(n5911) );
  DFFRX1 \CACHE_reg[2][58]  ( .D(n4672), .CK(clk), .RN(n516), .Q(
        \CACHE[2][58] ), .QN(n5912) );
  DFFRX1 \CACHE_reg[2][57]  ( .D(n4673), .CK(clk), .RN(n517), .Q(
        \CACHE[2][57] ), .QN(n5913) );
  DFFRX1 \CACHE_reg[2][56]  ( .D(n4674), .CK(clk), .RN(n517), .Q(
        \CACHE[2][56] ), .QN(n5914) );
  DFFRX1 \CACHE_reg[2][55]  ( .D(n4675), .CK(clk), .RN(n518), .Q(
        \CACHE[2][55] ), .QN(n5915) );
  DFFRX1 \CACHE_reg[2][54]  ( .D(n4676), .CK(clk), .RN(n519), .Q(
        \CACHE[2][54] ), .QN(n5916) );
  DFFRX1 \CACHE_reg[2][53]  ( .D(n4677), .CK(clk), .RN(n519), .Q(
        \CACHE[2][53] ), .QN(n5917) );
  DFFRX1 \CACHE_reg[2][52]  ( .D(n4678), .CK(clk), .RN(n520), .Q(
        \CACHE[2][52] ), .QN(n5918) );
  DFFRX1 \CACHE_reg[2][51]  ( .D(n4679), .CK(clk), .RN(n521), .Q(
        \CACHE[2][51] ), .QN(n5919) );
  DFFRX1 \CACHE_reg[2][50]  ( .D(n4680), .CK(clk), .RN(n521), .Q(
        \CACHE[2][50] ), .QN(n5920) );
  DFFRX1 \CACHE_reg[2][49]  ( .D(n4681), .CK(clk), .RN(n522), .Q(
        \CACHE[2][49] ), .QN(n5921) );
  DFFRX1 \CACHE_reg[2][48]  ( .D(n4682), .CK(clk), .RN(n523), .Q(
        \CACHE[2][48] ), .QN(n5922) );
  DFFRX1 \CACHE_reg[2][47]  ( .D(n4683), .CK(clk), .RN(n523), .Q(
        \CACHE[2][47] ), .QN(n5923) );
  DFFRX1 \CACHE_reg[2][46]  ( .D(n4684), .CK(clk), .RN(n524), .Q(
        \CACHE[2][46] ), .QN(n5924) );
  DFFRX1 \CACHE_reg[2][45]  ( .D(n4685), .CK(clk), .RN(n525), .Q(
        \CACHE[2][45] ), .QN(n5925) );
  DFFRX1 \CACHE_reg[2][44]  ( .D(n4686), .CK(clk), .RN(n525), .Q(
        \CACHE[2][44] ), .QN(n5926) );
  DFFRX1 \CACHE_reg[2][43]  ( .D(n4687), .CK(clk), .RN(n526), .Q(
        \CACHE[2][43] ), .QN(n5927) );
  DFFRX1 \CACHE_reg[2][42]  ( .D(n4688), .CK(clk), .RN(n527), .Q(
        \CACHE[2][42] ), .QN(n5928) );
  DFFRX1 \CACHE_reg[2][41]  ( .D(n4689), .CK(clk), .RN(n527), .Q(
        \CACHE[2][41] ), .QN(n5929) );
  DFFRX1 \CACHE_reg[2][40]  ( .D(n4690), .CK(clk), .RN(n528), .Q(
        \CACHE[2][40] ), .QN(n5930) );
  DFFRX1 \CACHE_reg[2][39]  ( .D(n4691), .CK(clk), .RN(n529), .Q(
        \CACHE[2][39] ), .QN(n5931) );
  DFFRX1 \CACHE_reg[2][38]  ( .D(n4692), .CK(clk), .RN(n529), .Q(
        \CACHE[2][38] ), .QN(n5932) );
  DFFRX1 \CACHE_reg[2][37]  ( .D(n4693), .CK(clk), .RN(n530), .Q(
        \CACHE[2][37] ), .QN(n5933) );
  DFFRX1 \CACHE_reg[2][36]  ( .D(n4694), .CK(clk), .RN(n531), .Q(
        \CACHE[2][36] ), .QN(n5934) );
  DFFRX1 \CACHE_reg[2][35]  ( .D(n4695), .CK(clk), .RN(n531), .Q(
        \CACHE[2][35] ), .QN(n5935) );
  DFFRX1 \CACHE_reg[2][34]  ( .D(n4696), .CK(clk), .RN(n532), .Q(
        \CACHE[2][34] ), .QN(n5936) );
  DFFRX1 \CACHE_reg[2][33]  ( .D(n4697), .CK(clk), .RN(n533), .Q(
        \CACHE[2][33] ), .QN(n5937) );
  DFFRX1 \CACHE_reg[2][32]  ( .D(n4698), .CK(clk), .RN(n533), .Q(
        \CACHE[2][32] ), .QN(n5938) );
  DFFRX1 \CACHE_reg[2][31]  ( .D(n4699), .CK(clk), .RN(n491), .Q(
        \CACHE[2][31] ), .QN(n5939) );
  DFFRX1 \CACHE_reg[2][30]  ( .D(n4700), .CK(clk), .RN(n3056), .Q(
        \CACHE[2][30] ), .QN(n5940) );
  DFFRX1 \CACHE_reg[2][29]  ( .D(n4701), .CK(clk), .RN(n493), .Q(
        \CACHE[2][29] ), .QN(n5941) );
  DFFRX1 \CACHE_reg[2][28]  ( .D(n4702), .CK(clk), .RN(n493), .Q(
        \CACHE[2][28] ), .QN(n5942) );
  DFFRX1 \CACHE_reg[2][27]  ( .D(n4703), .CK(clk), .RN(n494), .Q(
        \CACHE[2][27] ), .QN(n5943) );
  DFFRX1 \CACHE_reg[2][26]  ( .D(n4704), .CK(clk), .RN(n495), .Q(
        \CACHE[2][26] ), .QN(n5944) );
  DFFRX1 \CACHE_reg[2][25]  ( .D(n4705), .CK(clk), .RN(n495), .Q(
        \CACHE[2][25] ), .QN(n5945) );
  DFFRX1 \CACHE_reg[2][24]  ( .D(n4706), .CK(clk), .RN(n496), .Q(
        \CACHE[2][24] ), .QN(n5946) );
  DFFRX1 \CACHE_reg[2][23]  ( .D(n4707), .CK(clk), .RN(n497), .Q(
        \CACHE[2][23] ), .QN(n5947) );
  DFFRX1 \CACHE_reg[2][22]  ( .D(n4708), .CK(clk), .RN(n497), .Q(
        \CACHE[2][22] ), .QN(n5948) );
  DFFRX1 \CACHE_reg[2][21]  ( .D(n4709), .CK(clk), .RN(n498), .Q(
        \CACHE[2][21] ), .QN(n5949) );
  DFFRX1 \CACHE_reg[2][20]  ( .D(n4710), .CK(clk), .RN(n499), .Q(
        \CACHE[2][20] ), .QN(n5950) );
  DFFRX1 \CACHE_reg[2][19]  ( .D(n4711), .CK(clk), .RN(n499), .Q(
        \CACHE[2][19] ), .QN(n5951) );
  DFFRX1 \CACHE_reg[2][18]  ( .D(n4712), .CK(clk), .RN(n500), .Q(
        \CACHE[2][18] ), .QN(n5952) );
  DFFRX1 \CACHE_reg[2][17]  ( .D(n4713), .CK(clk), .RN(n501), .Q(
        \CACHE[2][17] ), .QN(n5953) );
  DFFRX1 \CACHE_reg[2][16]  ( .D(n4714), .CK(clk), .RN(n501), .Q(
        \CACHE[2][16] ), .QN(n5954) );
  DFFRX1 \CACHE_reg[2][15]  ( .D(n4715), .CK(clk), .RN(n502), .Q(
        \CACHE[2][15] ), .QN(n5955) );
  DFFRX1 \CACHE_reg[2][14]  ( .D(n4716), .CK(clk), .RN(n503), .Q(
        \CACHE[2][14] ), .QN(n5956) );
  DFFRX1 \CACHE_reg[2][13]  ( .D(n4717), .CK(clk), .RN(n503), .Q(
        \CACHE[2][13] ), .QN(n5957) );
  DFFRX1 \CACHE_reg[2][12]  ( .D(n4718), .CK(clk), .RN(n504), .Q(
        \CACHE[2][12] ), .QN(n5958) );
  DFFRX1 \CACHE_reg[2][11]  ( .D(n4719), .CK(clk), .RN(n505), .Q(
        \CACHE[2][11] ), .QN(n5959) );
  DFFRX1 \CACHE_reg[2][10]  ( .D(n4720), .CK(clk), .RN(n505), .Q(
        \CACHE[2][10] ), .QN(n5960) );
  DFFRX1 \CACHE_reg[2][9]  ( .D(n4721), .CK(clk), .RN(n506), .Q(\CACHE[2][9] ), 
        .QN(n5961) );
  DFFRX1 \CACHE_reg[2][8]  ( .D(n4722), .CK(clk), .RN(n507), .Q(\CACHE[2][8] ), 
        .QN(n5962) );
  DFFRX1 \CACHE_reg[2][7]  ( .D(n4723), .CK(clk), .RN(n507), .Q(\CACHE[2][7] ), 
        .QN(n5963) );
  DFFRX1 \CACHE_reg[2][6]  ( .D(n4724), .CK(clk), .RN(n508), .Q(\CACHE[2][6] ), 
        .QN(n5964) );
  DFFRX1 \CACHE_reg[2][5]  ( .D(n4725), .CK(clk), .RN(n509), .Q(\CACHE[2][5] ), 
        .QN(n5965) );
  DFFRX1 \CACHE_reg[2][4]  ( .D(n4726), .CK(clk), .RN(n509), .Q(\CACHE[2][4] ), 
        .QN(n5966) );
  DFFRX1 \CACHE_reg[2][3]  ( .D(n4727), .CK(clk), .RN(n510), .Q(\CACHE[2][3] ), 
        .QN(n5967) );
  DFFRX1 \CACHE_reg[2][2]  ( .D(n4728), .CK(clk), .RN(n511), .Q(\CACHE[2][2] ), 
        .QN(n5968) );
  DFFRX1 \CACHE_reg[2][1]  ( .D(n4729), .CK(clk), .RN(n511), .Q(\CACHE[2][1] ), 
        .QN(n5969) );
  DFFRX1 \CACHE_reg[2][0]  ( .D(n4730), .CK(clk), .RN(n512), .Q(\CACHE[2][0] ), 
        .QN(n5970) );
  AND2X2 U3 ( .A(n3764), .B(mem_ready), .Y(n3741) );
  OR2X1 U4 ( .A(n3765), .B(n473), .Y(n1) );
  OR2X1 U5 ( .A(n3569), .B(n399), .Y(n2) );
  OR2X1 U6 ( .A(n3514), .B(n402), .Y(n3) );
  OR2X1 U7 ( .A(n3459), .B(n403), .Y(n4) );
  OR2X1 U8 ( .A(n3444), .B(n404), .Y(n5) );
  OR2X1 U9 ( .A(n3439), .B(n405), .Y(n6) );
  OR2X1 U10 ( .A(n3434), .B(n405), .Y(n7) );
  OR2X1 U11 ( .A(n3429), .B(n406), .Y(n8) );
  OR2X1 U12 ( .A(n3424), .B(n407), .Y(n9) );
  OR2X1 U13 ( .A(n3419), .B(n408), .Y(n10) );
  OR2X1 U14 ( .A(n3413), .B(n409), .Y(n11) );
  OR2X1 U15 ( .A(n3564), .B(n399), .Y(n12) );
  OR2X1 U16 ( .A(n3559), .B(n400), .Y(n13) );
  OR2X1 U17 ( .A(n3554), .B(n401), .Y(n14) );
  OR2X1 U18 ( .A(n3549), .B(n401), .Y(n15) );
  OR2X1 U19 ( .A(n3544), .B(n401), .Y(n16) );
  OR2X1 U20 ( .A(n3539), .B(n401), .Y(n17) );
  OR2X1 U21 ( .A(n3534), .B(n401), .Y(n18) );
  OR2X1 U22 ( .A(n3529), .B(n402), .Y(n19) );
  OR2X1 U23 ( .A(n3524), .B(n402), .Y(n20) );
  OR2X1 U24 ( .A(n3519), .B(n402), .Y(n21) );
  OR2X1 U25 ( .A(n3509), .B(n402), .Y(n22) );
  OR2X1 U26 ( .A(n3504), .B(n402), .Y(n23) );
  OR2X1 U27 ( .A(n3499), .B(n402), .Y(n24) );
  OR2X1 U28 ( .A(n3494), .B(n402), .Y(n25) );
  OR2X1 U29 ( .A(n3489), .B(n402), .Y(n26) );
  OR2X1 U30 ( .A(n3484), .B(n402), .Y(n27) );
  OR2X1 U31 ( .A(n3479), .B(n402), .Y(n28) );
  OR2X1 U32 ( .A(n3474), .B(n402), .Y(n29) );
  OR2X1 U33 ( .A(n3469), .B(n403), .Y(n30) );
  OR2X1 U34 ( .A(n3464), .B(n403), .Y(n31) );
  OR2X1 U35 ( .A(n3454), .B(n403), .Y(n32) );
  OR2X1 U36 ( .A(n3449), .B(n403), .Y(n33) );
  OR2X1 U37 ( .A(n3567), .B(n403), .Y(n34) );
  OR2X1 U38 ( .A(n3512), .B(n403), .Y(n35) );
  OR2X1 U39 ( .A(n3457), .B(n403), .Y(n36) );
  OR2X1 U40 ( .A(n3442), .B(n403), .Y(n37) );
  OR2X1 U41 ( .A(n3437), .B(n403), .Y(n38) );
  OR2X1 U42 ( .A(n3432), .B(n403), .Y(n39) );
  OR2X1 U43 ( .A(n3427), .B(n403), .Y(n40) );
  OR2X1 U44 ( .A(n3422), .B(n404), .Y(n41) );
  OR2X1 U45 ( .A(n3417), .B(n404), .Y(n42) );
  OR2X1 U46 ( .A(n3410), .B(n404), .Y(n43) );
  OR2X1 U47 ( .A(n3562), .B(n404), .Y(n44) );
  OR2X1 U48 ( .A(n3557), .B(n404), .Y(n45) );
  OR2X1 U49 ( .A(n3552), .B(n404), .Y(n46) );
  OR2X1 U50 ( .A(n3547), .B(n404), .Y(n47) );
  OR2X1 U51 ( .A(n3542), .B(n404), .Y(n48) );
  OR2X1 U52 ( .A(n3537), .B(n404), .Y(n49) );
  OR2X1 U53 ( .A(n3532), .B(n404), .Y(n50) );
  OR2X1 U54 ( .A(n3527), .B(n404), .Y(n51) );
  OR2X1 U55 ( .A(n3522), .B(n405), .Y(n52) );
  OR2X1 U56 ( .A(n3517), .B(n405), .Y(n53) );
  OR2X1 U57 ( .A(n3507), .B(n405), .Y(n54) );
  OR2X1 U58 ( .A(n3502), .B(n405), .Y(n55) );
  OR2X1 U59 ( .A(n3497), .B(n405), .Y(n56) );
  OR2X1 U60 ( .A(n3492), .B(n405), .Y(n57) );
  OR2X1 U61 ( .A(n3487), .B(n405), .Y(n58) );
  OR2X1 U62 ( .A(n3482), .B(n405), .Y(n59) );
  OR2X1 U63 ( .A(n3477), .B(n405), .Y(n60) );
  OR2X1 U64 ( .A(n3472), .B(n405), .Y(n61) );
  OR2X1 U65 ( .A(n3467), .B(n406), .Y(n62) );
  OR2X1 U66 ( .A(n3462), .B(n406), .Y(n63) );
  OR2X1 U67 ( .A(n3452), .B(n406), .Y(n64) );
  OR2X1 U68 ( .A(n3447), .B(n406), .Y(n65) );
  OR2X1 U69 ( .A(n3566), .B(n406), .Y(n66) );
  OR2X1 U70 ( .A(n3511), .B(n406), .Y(n67) );
  OR2X1 U71 ( .A(n3456), .B(n406), .Y(n68) );
  OR2X1 U72 ( .A(n3441), .B(n406), .Y(n69) );
  OR2X1 U73 ( .A(n3436), .B(n406), .Y(n70) );
  OR2X1 U74 ( .A(n3431), .B(n406), .Y(n71) );
  OR2X1 U75 ( .A(n3426), .B(n406), .Y(n72) );
  OR2X1 U76 ( .A(n3421), .B(n407), .Y(n73) );
  OR2X1 U77 ( .A(n3416), .B(n407), .Y(n74) );
  OR2X1 U78 ( .A(n3408), .B(n407), .Y(n75) );
  OR2X1 U79 ( .A(n3561), .B(n407), .Y(n76) );
  OR2X1 U80 ( .A(n3556), .B(n407), .Y(n77) );
  OR2X1 U81 ( .A(n3551), .B(n407), .Y(n78) );
  OR2X1 U82 ( .A(n3546), .B(n407), .Y(n79) );
  OR2X1 U83 ( .A(n3541), .B(n407), .Y(n80) );
  OR2X1 U84 ( .A(n3536), .B(n407), .Y(n81) );
  OR2X1 U85 ( .A(n3531), .B(n407), .Y(n82) );
  OR2X1 U86 ( .A(n3526), .B(n407), .Y(n83) );
  OR2X1 U87 ( .A(n3521), .B(n408), .Y(n84) );
  OR2X1 U88 ( .A(n3516), .B(n408), .Y(n85) );
  OR2X1 U89 ( .A(n3506), .B(n408), .Y(n86) );
  OR2X1 U90 ( .A(n3501), .B(n408), .Y(n87) );
  OR2X1 U91 ( .A(n3496), .B(n408), .Y(n88) );
  OR2X1 U92 ( .A(n3491), .B(n408), .Y(n89) );
  OR2X1 U93 ( .A(n3486), .B(n408), .Y(n90) );
  OR2X1 U94 ( .A(n3481), .B(n408), .Y(n91) );
  OR2X1 U95 ( .A(n3476), .B(n408), .Y(n92) );
  OR2X1 U96 ( .A(n3471), .B(n408), .Y(n93) );
  OR2X1 U97 ( .A(n3466), .B(n408), .Y(n94) );
  OR2X1 U98 ( .A(n3461), .B(n409), .Y(n95) );
  OR2X1 U99 ( .A(n3451), .B(n409), .Y(n96) );
  OR2X1 U100 ( .A(n3446), .B(n409), .Y(n97) );
  OR2X1 U101 ( .A(n3570), .B(n409), .Y(n98) );
  OR2X1 U102 ( .A(n3515), .B(n409), .Y(n99) );
  OR2X1 U103 ( .A(n3460), .B(n409), .Y(n100) );
  OR2X1 U104 ( .A(n3445), .B(n409), .Y(n101) );
  OR2X1 U105 ( .A(n3440), .B(n399), .Y(n102) );
  OR2X1 U106 ( .A(n3435), .B(n399), .Y(n103) );
  OR2X1 U107 ( .A(n3430), .B(n399), .Y(n104) );
  OR2X1 U108 ( .A(n3425), .B(n399), .Y(n105) );
  OR2X1 U109 ( .A(n3420), .B(n399), .Y(n106) );
  OR2X1 U110 ( .A(n3415), .B(n399), .Y(n107) );
  OR2X1 U111 ( .A(n3565), .B(n399), .Y(n108) );
  OR2X1 U112 ( .A(n3560), .B(n399), .Y(n109) );
  OR2X1 U113 ( .A(n3555), .B(n399), .Y(n110) );
  OR2X1 U114 ( .A(n3550), .B(n399), .Y(n111) );
  OR2X1 U115 ( .A(n3545), .B(n400), .Y(n112) );
  OR2X1 U116 ( .A(n3540), .B(n400), .Y(n113) );
  OR2X1 U117 ( .A(n3535), .B(n400), .Y(n114) );
  OR2X1 U118 ( .A(n3530), .B(n400), .Y(n115) );
  OR2X1 U119 ( .A(n3525), .B(n400), .Y(n116) );
  OR2X1 U120 ( .A(n3520), .B(n400), .Y(n117) );
  OR2X1 U121 ( .A(n3510), .B(n400), .Y(n118) );
  OR2X1 U122 ( .A(n3505), .B(n400), .Y(n119) );
  OR2X1 U123 ( .A(n3500), .B(n400), .Y(n120) );
  OR2X1 U124 ( .A(n3495), .B(n400), .Y(n121) );
  OR2X1 U125 ( .A(n3490), .B(n400), .Y(n122) );
  OR2X1 U126 ( .A(n3485), .B(n401), .Y(n123) );
  OR2X1 U127 ( .A(n3480), .B(n401), .Y(n124) );
  OR2X1 U128 ( .A(n3475), .B(n401), .Y(n125) );
  OR2X1 U129 ( .A(n3470), .B(n401), .Y(n126) );
  OR2X1 U130 ( .A(n3465), .B(n401), .Y(n127) );
  OR2X1 U131 ( .A(n3455), .B(n401), .Y(n128) );
  OR2X1 U132 ( .A(n3450), .B(n401), .Y(n129) );
  OR2X1 U133 ( .A(n3765), .B(n435), .Y(n130) );
  OR2X1 U134 ( .A(n3765), .B(n460), .Y(n131) );
  AOI22X1 U135 ( .A0(N59), .A1(n412), .B0(proc_addr[5]), .B1(mem_read), .Y(
        n132) );
  AOI22X1 U136 ( .A0(N58), .A1(n412), .B0(proc_addr[6]), .B1(mem_read), .Y(
        n133) );
  AOI22X1 U137 ( .A0(N57), .A1(n412), .B0(proc_addr[7]), .B1(mem_read), .Y(
        n134) );
  AOI22X1 U138 ( .A0(N56), .A1(n315), .B0(proc_addr[8]), .B1(mem_read), .Y(
        n135) );
  AOI22X1 U139 ( .A0(N55), .A1(mem_write), .B0(proc_addr[9]), .B1(mem_read), 
        .Y(n136) );
  AOI22X1 U140 ( .A0(N54), .A1(n410), .B0(proc_addr[10]), .B1(mem_read), .Y(
        n137) );
  AOI22X1 U141 ( .A0(N53), .A1(n414), .B0(proc_addr[11]), .B1(mem_read), .Y(
        n138) );
  AOI22X1 U142 ( .A0(N52), .A1(n410), .B0(proc_addr[12]), .B1(mem_read), .Y(
        n139) );
  AOI22X1 U143 ( .A0(N51), .A1(n414), .B0(proc_addr[13]), .B1(mem_read), .Y(
        n140) );
  AOI22X1 U144 ( .A0(N50), .A1(n315), .B0(proc_addr[14]), .B1(mem_read), .Y(
        n141) );
  AOI22X1 U145 ( .A0(N49), .A1(n410), .B0(proc_addr[15]), .B1(mem_read), .Y(
        n142) );
  AOI22X1 U146 ( .A0(N48), .A1(n410), .B0(proc_addr[16]), .B1(mem_read), .Y(
        n143) );
  AOI22X1 U147 ( .A0(N47), .A1(n410), .B0(proc_addr[17]), .B1(mem_read), .Y(
        n144) );
  AOI22X1 U148 ( .A0(N46), .A1(mem_write), .B0(proc_addr[18]), .B1(mem_read), 
        .Y(n145) );
  AOI22X1 U149 ( .A0(N45), .A1(mem_write), .B0(proc_addr[19]), .B1(mem_read), 
        .Y(n146) );
  AOI22X1 U150 ( .A0(N44), .A1(n414), .B0(proc_addr[20]), .B1(mem_read), .Y(
        n147) );
  AOI22X1 U151 ( .A0(N43), .A1(n413), .B0(proc_addr[21]), .B1(mem_read), .Y(
        n148) );
  AOI22X1 U152 ( .A0(N42), .A1(mem_write), .B0(proc_addr[22]), .B1(mem_read), 
        .Y(n149) );
  AOI22X1 U153 ( .A0(N41), .A1(mem_write), .B0(proc_addr[23]), .B1(mem_read), 
        .Y(n150) );
  AOI22X1 U154 ( .A0(N40), .A1(mem_write), .B0(proc_addr[24]), .B1(mem_read), 
        .Y(n151) );
  AOI22X1 U155 ( .A0(N39), .A1(n412), .B0(proc_addr[25]), .B1(mem_read), .Y(
        n152) );
  AOI22X1 U156 ( .A0(N38), .A1(n412), .B0(proc_addr[26]), .B1(mem_read), .Y(
        n153) );
  AOI22X1 U157 ( .A0(N37), .A1(n412), .B0(proc_addr[27]), .B1(mem_read), .Y(
        n154) );
  AOI22X1 U158 ( .A0(N36), .A1(n412), .B0(proc_addr[28]), .B1(mem_read), .Y(
        n155) );
  AOI22X1 U159 ( .A0(N35), .A1(n412), .B0(proc_addr[29]), .B1(mem_read), .Y(
        n156) );
  AOI22X2 U160 ( .A0(proc_addr[29]), .A1(n391), .B0(n3742), .B1(N35), .Y(n3577) );
  AOI22X2 U161 ( .A0(proc_addr[28]), .A1(n391), .B0(n3742), .B1(N36), .Y(n3578) );
  AOI22X2 U162 ( .A0(proc_addr[27]), .A1(n391), .B0(n3742), .B1(N37), .Y(n3579) );
  AOI22X2 U163 ( .A0(proc_addr[26]), .A1(n391), .B0(n3742), .B1(N38), .Y(n3580) );
  AOI22X2 U164 ( .A0(proc_addr[25]), .A1(n391), .B0(n3742), .B1(N39), .Y(n3581) );
  AOI22X2 U165 ( .A0(proc_addr[24]), .A1(n391), .B0(n3742), .B1(N40), .Y(n3582) );
  AOI22X2 U166 ( .A0(proc_addr[23]), .A1(n391), .B0(n3742), .B1(N41), .Y(n3583) );
  AOI22X2 U167 ( .A0(proc_addr[22]), .A1(n391), .B0(n3742), .B1(N42), .Y(n3584) );
  AOI22X2 U168 ( .A0(proc_addr[21]), .A1(n391), .B0(n3742), .B1(N43), .Y(n3585) );
  AOI22X2 U169 ( .A0(proc_addr[20]), .A1(n391), .B0(n3742), .B1(N44), .Y(n3586) );
  CLKBUFX3 U170 ( .A(n3741), .Y(n391) );
  AOI22X2 U171 ( .A0(proc_addr[19]), .A1(n391), .B0(n3742), .B1(N45), .Y(n3587) );
  AOI22X2 U172 ( .A0(proc_addr[18]), .A1(n391), .B0(n3742), .B1(N46), .Y(n3588) );
  AOI22X2 U173 ( .A0(proc_addr[17]), .A1(n392), .B0(n3742), .B1(N47), .Y(n3589) );
  AOI22X2 U174 ( .A0(proc_addr[16]), .A1(n392), .B0(n3742), .B1(N48), .Y(n3590) );
  AOI22X2 U175 ( .A0(proc_addr[15]), .A1(n392), .B0(n3742), .B1(N49), .Y(n3591) );
  AOI22X2 U176 ( .A0(proc_addr[14]), .A1(n392), .B0(n3742), .B1(N50), .Y(n3592) );
  AOI22X2 U177 ( .A0(proc_addr[13]), .A1(n392), .B0(n3742), .B1(N51), .Y(n3593) );
  AOI22X2 U178 ( .A0(proc_addr[12]), .A1(n392), .B0(n3742), .B1(N52), .Y(n3594) );
  AOI22X2 U179 ( .A0(proc_addr[11]), .A1(n392), .B0(n3742), .B1(N53), .Y(n3595) );
  AOI222X4 U180 ( .A0(mem_rdata[127]), .A1(n397), .B0(n3745), .B1(N60), .C0(
        proc_wdata[31]), .C1(n3746), .Y(n3602) );
  AOI222X4 U181 ( .A0(mem_rdata[126]), .A1(n396), .B0(n3745), .B1(N61), .C0(
        proc_wdata[30]), .C1(n3746), .Y(n3603) );
  AOI222X4 U182 ( .A0(mem_rdata[125]), .A1(n394), .B0(n3745), .B1(N62), .C0(
        proc_wdata[29]), .C1(n3746), .Y(n3604) );
  AOI222X4 U183 ( .A0(mem_rdata[124]), .A1(n3741), .B0(n3745), .B1(N63), .C0(
        proc_wdata[28]), .C1(n3746), .Y(n3605) );
  AOI222X4 U184 ( .A0(mem_rdata[123]), .A1(n397), .B0(n3745), .B1(N64), .C0(
        proc_wdata[27]), .C1(n3746), .Y(n3606) );
  AOI222X4 U185 ( .A0(mem_rdata[122]), .A1(n396), .B0(n3745), .B1(N65), .C0(
        proc_wdata[26]), .C1(n3746), .Y(n3607) );
  AOI222X4 U186 ( .A0(mem_rdata[121]), .A1(n394), .B0(n3745), .B1(N66), .C0(
        proc_wdata[25]), .C1(n3746), .Y(n3608) );
  AOI222X4 U187 ( .A0(mem_rdata[120]), .A1(n394), .B0(n3745), .B1(N67), .C0(
        proc_wdata[24]), .C1(n3746), .Y(n3609) );
  AOI222X4 U188 ( .A0(mem_rdata[119]), .A1(n398), .B0(n3745), .B1(N68), .C0(
        proc_wdata[23]), .C1(n3746), .Y(n3610) );
  AOI222X4 U189 ( .A0(mem_rdata[118]), .A1(n397), .B0(n3745), .B1(N69), .C0(
        proc_wdata[22]), .C1(n3746), .Y(n3611) );
  AOI222X4 U190 ( .A0(mem_rdata[117]), .A1(n393), .B0(n3745), .B1(N70), .C0(
        proc_wdata[21]), .C1(n3746), .Y(n3612) );
  AOI222X4 U191 ( .A0(mem_rdata[116]), .A1(n396), .B0(n3745), .B1(N71), .C0(
        proc_wdata[20]), .C1(n3746), .Y(n3613) );
  AOI222X4 U192 ( .A0(mem_rdata[115]), .A1(n392), .B0(n3745), .B1(N72), .C0(
        proc_wdata[19]), .C1(n3746), .Y(n3614) );
  AOI222X4 U193 ( .A0(mem_rdata[114]), .A1(n391), .B0(n3745), .B1(N73), .C0(
        proc_wdata[18]), .C1(n3746), .Y(n3615) );
  AOI222X4 U194 ( .A0(mem_rdata[113]), .A1(n395), .B0(n3745), .B1(N74), .C0(
        proc_wdata[17]), .C1(n3746), .Y(n3616) );
  AOI222X4 U195 ( .A0(mem_rdata[112]), .A1(n397), .B0(n3745), .B1(N75), .C0(
        proc_wdata[16]), .C1(n3746), .Y(n3617) );
  AOI222X4 U196 ( .A0(mem_rdata[111]), .A1(n393), .B0(n3745), .B1(N76), .C0(
        proc_wdata[15]), .C1(n3746), .Y(n3618) );
  AOI222X4 U197 ( .A0(mem_rdata[110]), .A1(n396), .B0(n3745), .B1(N77), .C0(
        proc_wdata[14]), .C1(n3746), .Y(n3619) );
  AOI222X4 U198 ( .A0(mem_rdata[109]), .A1(n392), .B0(n3745), .B1(N78), .C0(
        proc_wdata[13]), .C1(n3746), .Y(n3620) );
  AOI222X4 U199 ( .A0(mem_rdata[108]), .A1(n391), .B0(n3745), .B1(N79), .C0(
        proc_wdata[12]), .C1(n3746), .Y(n3621) );
  AOI222X4 U200 ( .A0(mem_rdata[107]), .A1(n3741), .B0(n3745), .B1(N80), .C0(
        proc_wdata[11]), .C1(n3746), .Y(n3622) );
  AOI222X4 U201 ( .A0(mem_rdata[106]), .A1(n3741), .B0(n3745), .B1(N81), .C0(
        proc_wdata[10]), .C1(n3746), .Y(n3623) );
  AOI222X4 U202 ( .A0(mem_rdata[105]), .A1(n3741), .B0(n3745), .B1(N82), .C0(
        proc_wdata[9]), .C1(n3746), .Y(n3624) );
  AOI222X4 U203 ( .A0(mem_rdata[104]), .A1(n3741), .B0(n3745), .B1(N83), .C0(
        proc_wdata[8]), .C1(n3746), .Y(n3625) );
  AOI222X4 U204 ( .A0(mem_rdata[103]), .A1(n3741), .B0(n3745), .B1(N84), .C0(
        proc_wdata[7]), .C1(n3746), .Y(n3626) );
  AOI222X4 U205 ( .A0(mem_rdata[102]), .A1(n392), .B0(n3745), .B1(N85), .C0(
        proc_wdata[6]), .C1(n3746), .Y(n3627) );
  AOI222X4 U206 ( .A0(mem_rdata[101]), .A1(n391), .B0(n3745), .B1(N86), .C0(
        proc_wdata[5]), .C1(n3746), .Y(n3628) );
  AOI222X4 U207 ( .A0(mem_rdata[100]), .A1(n398), .B0(n3745), .B1(N87), .C0(
        proc_wdata[4]), .C1(n3746), .Y(n3629) );
  AOI222X4 U208 ( .A0(mem_rdata[99]), .A1(n395), .B0(n3745), .B1(N88), .C0(
        proc_wdata[3]), .C1(n3746), .Y(n3630) );
  AOI222X4 U209 ( .A0(mem_rdata[98]), .A1(n397), .B0(n3745), .B1(N89), .C0(
        proc_wdata[2]), .C1(n3746), .Y(n3631) );
  AOI222X4 U210 ( .A0(mem_rdata[97]), .A1(n393), .B0(n3745), .B1(N90), .C0(
        proc_wdata[1]), .C1(n3746), .Y(n3632) );
  AOI222X4 U211 ( .A0(mem_rdata[96]), .A1(n393), .B0(n3745), .B1(N91), .C0(
        proc_wdata[0]), .C1(n3746), .Y(n3633) );
  AOI222X4 U212 ( .A0(n398), .A1(mem_rdata[95]), .B0(proc_wdata[31]), .B1(
        n3750), .C0(N92), .C1(n3751), .Y(n3634) );
  AOI222X4 U213 ( .A0(n398), .A1(mem_rdata[94]), .B0(proc_wdata[30]), .B1(
        n3750), .C0(N93), .C1(n3751), .Y(n3635) );
  AOI222X4 U214 ( .A0(n398), .A1(mem_rdata[93]), .B0(proc_wdata[29]), .B1(
        n3750), .C0(N94), .C1(n3751), .Y(n3636) );
  AOI222X4 U215 ( .A0(n398), .A1(mem_rdata[92]), .B0(proc_wdata[28]), .B1(
        n3750), .C0(N95), .C1(n3751), .Y(n3637) );
  AOI222X4 U216 ( .A0(n398), .A1(mem_rdata[91]), .B0(proc_wdata[27]), .B1(
        n3750), .C0(N96), .C1(n3751), .Y(n3638) );
  AOI222X4 U217 ( .A0(n397), .A1(mem_rdata[90]), .B0(proc_wdata[26]), .B1(
        n3750), .C0(N97), .C1(n3751), .Y(n3639) );
  AOI222X4 U218 ( .A0(n398), .A1(mem_rdata[89]), .B0(proc_wdata[25]), .B1(
        n3750), .C0(N98), .C1(n3751), .Y(n3640) );
  AOI222X4 U219 ( .A0(n3741), .A1(mem_rdata[88]), .B0(proc_wdata[24]), .B1(
        n3750), .C0(N99), .C1(n3751), .Y(n3641) );
  AOI222X4 U220 ( .A0(n397), .A1(mem_rdata[87]), .B0(proc_wdata[23]), .B1(
        n3750), .C0(N100), .C1(n3751), .Y(n3642) );
  AOI222X4 U221 ( .A0(n398), .A1(mem_rdata[86]), .B0(proc_wdata[22]), .B1(
        n3750), .C0(N101), .C1(n3751), .Y(n3643) );
  AOI222X4 U222 ( .A0(n397), .A1(mem_rdata[85]), .B0(proc_wdata[21]), .B1(
        n3750), .C0(N102), .C1(n3751), .Y(n3644) );
  AOI222X4 U223 ( .A0(n397), .A1(mem_rdata[84]), .B0(proc_wdata[20]), .B1(
        n3750), .C0(N103), .C1(n3751), .Y(n3645) );
  AOI222X4 U224 ( .A0(n398), .A1(mem_rdata[83]), .B0(proc_wdata[19]), .B1(
        n3750), .C0(N104), .C1(n3751), .Y(n3646) );
  AOI222X4 U225 ( .A0(n397), .A1(mem_rdata[82]), .B0(proc_wdata[18]), .B1(
        n3750), .C0(N105), .C1(n3751), .Y(n3647) );
  AOI222X4 U226 ( .A0(n397), .A1(mem_rdata[81]), .B0(proc_wdata[17]), .B1(
        n3750), .C0(N106), .C1(n3751), .Y(n3648) );
  AOI222X4 U227 ( .A0(n3741), .A1(mem_rdata[80]), .B0(proc_wdata[16]), .B1(
        n3750), .C0(N107), .C1(n3751), .Y(n3649) );
  AOI222X4 U228 ( .A0(n397), .A1(mem_rdata[79]), .B0(proc_wdata[15]), .B1(
        n3750), .C0(N108), .C1(n3751), .Y(n3650) );
  AOI222X4 U229 ( .A0(n397), .A1(mem_rdata[78]), .B0(proc_wdata[14]), .B1(
        n3750), .C0(N109), .C1(n3751), .Y(n3651) );
  AOI222X4 U230 ( .A0(n398), .A1(mem_rdata[77]), .B0(proc_wdata[13]), .B1(
        n3750), .C0(N110), .C1(n3751), .Y(n3652) );
  AOI222X4 U231 ( .A0(n397), .A1(mem_rdata[76]), .B0(proc_wdata[12]), .B1(
        n3750), .C0(N111), .C1(n3751), .Y(n3653) );
  AOI222X4 U232 ( .A0(n397), .A1(mem_rdata[75]), .B0(proc_wdata[11]), .B1(
        n3750), .C0(N112), .C1(n3751), .Y(n3654) );
  AOI222X4 U233 ( .A0(n398), .A1(mem_rdata[74]), .B0(proc_wdata[10]), .B1(
        n3750), .C0(N113), .C1(n3751), .Y(n3655) );
  AOI222X4 U234 ( .A0(n397), .A1(mem_rdata[73]), .B0(proc_wdata[9]), .B1(n3750), .C0(N114), .C1(n3751), .Y(n3656) );
  AOI222X4 U235 ( .A0(n398), .A1(mem_rdata[72]), .B0(proc_wdata[8]), .B1(n3750), .C0(N115), .C1(n3751), .Y(n3657) );
  AOI222X4 U236 ( .A0(n398), .A1(mem_rdata[71]), .B0(proc_wdata[7]), .B1(n3750), .C0(N116), .C1(n3751), .Y(n3658) );
  AOI222X4 U237 ( .A0(n395), .A1(mem_rdata[70]), .B0(proc_wdata[6]), .B1(n3750), .C0(N117), .C1(n3751), .Y(n3659) );
  AOI222X4 U238 ( .A0(n397), .A1(mem_rdata[69]), .B0(proc_wdata[5]), .B1(n3750), .C0(N118), .C1(n3751), .Y(n3660) );
  AOI222X4 U239 ( .A0(n398), .A1(mem_rdata[68]), .B0(proc_wdata[4]), .B1(n3750), .C0(N119), .C1(n3751), .Y(n3661) );
  AOI222X4 U240 ( .A0(n397), .A1(mem_rdata[67]), .B0(proc_wdata[3]), .B1(n3750), .C0(N120), .C1(n3751), .Y(n3662) );
  AOI222X4 U241 ( .A0(n397), .A1(mem_rdata[66]), .B0(proc_wdata[2]), .B1(n3750), .C0(N121), .C1(n3751), .Y(n3663) );
  AOI222X4 U242 ( .A0(n398), .A1(mem_rdata[65]), .B0(proc_wdata[1]), .B1(n3750), .C0(N122), .C1(n3751), .Y(n3664) );
  AOI222X4 U243 ( .A0(n393), .A1(mem_rdata[64]), .B0(proc_wdata[0]), .B1(n3750), .C0(N123), .C1(n3751), .Y(n3665) );
  AOI222X4 U244 ( .A0(mem_rdata[63]), .A1(n396), .B0(n3753), .B1(N124), .C0(
        n3754), .C1(proc_wdata[31]), .Y(n3666) );
  AOI222X4 U245 ( .A0(mem_rdata[62]), .A1(n394), .B0(n3753), .B1(N125), .C0(
        n3754), .C1(proc_wdata[30]), .Y(n3667) );
  AOI222X4 U246 ( .A0(mem_rdata[61]), .A1(n392), .B0(n3753), .B1(N126), .C0(
        n3754), .C1(proc_wdata[29]), .Y(n3668) );
  AOI222X4 U247 ( .A0(mem_rdata[60]), .A1(n391), .B0(n3753), .B1(N127), .C0(
        n3754), .C1(proc_wdata[28]), .Y(n3669) );
  AOI222X4 U248 ( .A0(mem_rdata[59]), .A1(n398), .B0(n3753), .B1(N128), .C0(
        n3754), .C1(proc_wdata[27]), .Y(n3670) );
  AOI222X4 U249 ( .A0(mem_rdata[58]), .A1(n393), .B0(n3753), .B1(N129), .C0(
        n3754), .C1(proc_wdata[26]), .Y(n3671) );
  AOI222X4 U250 ( .A0(mem_rdata[57]), .A1(n394), .B0(n3753), .B1(N130), .C0(
        n3754), .C1(proc_wdata[25]), .Y(n3672) );
  AOI222X4 U251 ( .A0(mem_rdata[56]), .A1(n395), .B0(n3753), .B1(N131), .C0(
        n3754), .C1(proc_wdata[24]), .Y(n3673) );
  AOI222X4 U252 ( .A0(mem_rdata[55]), .A1(n394), .B0(n3753), .B1(N132), .C0(
        n3754), .C1(proc_wdata[23]), .Y(n3674) );
  AOI222X4 U253 ( .A0(mem_rdata[54]), .A1(n394), .B0(n3753), .B1(N133), .C0(
        n3754), .C1(proc_wdata[22]), .Y(n3675) );
  AOI222X4 U254 ( .A0(mem_rdata[53]), .A1(n393), .B0(n3753), .B1(N134), .C0(
        n3754), .C1(proc_wdata[21]), .Y(n3676) );
  AOI222X4 U255 ( .A0(mem_rdata[52]), .A1(n394), .B0(n3753), .B1(N135), .C0(
        n3754), .C1(proc_wdata[20]), .Y(n3677) );
  AOI222X4 U256 ( .A0(mem_rdata[51]), .A1(n394), .B0(n3753), .B1(N136), .C0(
        n3754), .C1(proc_wdata[19]), .Y(n3678) );
  AOI222X4 U257 ( .A0(mem_rdata[50]), .A1(n393), .B0(n3753), .B1(N137), .C0(
        n3754), .C1(proc_wdata[18]), .Y(n3679) );
  AOI222X4 U258 ( .A0(mem_rdata[49]), .A1(n394), .B0(n3753), .B1(N138), .C0(
        n3754), .C1(proc_wdata[17]), .Y(n3680) );
  AOI222X4 U259 ( .A0(mem_rdata[48]), .A1(n394), .B0(n3753), .B1(N139), .C0(
        n3754), .C1(proc_wdata[16]), .Y(n3681) );
  AOI222X4 U260 ( .A0(mem_rdata[47]), .A1(n393), .B0(n3753), .B1(N140), .C0(
        n3754), .C1(proc_wdata[15]), .Y(n3682) );
  AOI222X4 U261 ( .A0(mem_rdata[46]), .A1(n394), .B0(n3753), .B1(N141), .C0(
        n3754), .C1(proc_wdata[14]), .Y(n3683) );
  AOI222X4 U262 ( .A0(mem_rdata[45]), .A1(n394), .B0(n3753), .B1(N142), .C0(
        n3754), .C1(proc_wdata[13]), .Y(n3684) );
  AOI222X4 U263 ( .A0(mem_rdata[44]), .A1(n393), .B0(n3753), .B1(N143), .C0(
        n3754), .C1(proc_wdata[12]), .Y(n3685) );
  AOI222X4 U264 ( .A0(mem_rdata[43]), .A1(n393), .B0(n3753), .B1(N144), .C0(
        n3754), .C1(proc_wdata[11]), .Y(n3686) );
  AOI222X4 U265 ( .A0(mem_rdata[42]), .A1(n393), .B0(n3753), .B1(N145), .C0(
        n3754), .C1(proc_wdata[10]), .Y(n3687) );
  AOI222X4 U266 ( .A0(mem_rdata[41]), .A1(n393), .B0(n3753), .B1(N146), .C0(
        n3754), .C1(proc_wdata[9]), .Y(n3688) );
  AOI222X4 U267 ( .A0(mem_rdata[40]), .A1(n395), .B0(n3753), .B1(N147), .C0(
        n3754), .C1(proc_wdata[8]), .Y(n3689) );
  AOI222X4 U268 ( .A0(mem_rdata[39]), .A1(n395), .B0(n3753), .B1(N148), .C0(
        n3754), .C1(proc_wdata[7]), .Y(n3690) );
  AOI222X4 U269 ( .A0(mem_rdata[38]), .A1(n393), .B0(n3753), .B1(N149), .C0(
        n3754), .C1(proc_wdata[6]), .Y(n3691) );
  AOI222X4 U270 ( .A0(mem_rdata[37]), .A1(n395), .B0(n3753), .B1(N150), .C0(
        n3754), .C1(proc_wdata[5]), .Y(n3692) );
  AOI222X4 U271 ( .A0(mem_rdata[36]), .A1(n395), .B0(n3753), .B1(N151), .C0(
        n3754), .C1(proc_wdata[4]), .Y(n3693) );
  AOI222X4 U272 ( .A0(mem_rdata[35]), .A1(n393), .B0(n3753), .B1(N152), .C0(
        n3754), .C1(proc_wdata[3]), .Y(n3694) );
  AOI222X4 U273 ( .A0(mem_rdata[34]), .A1(n394), .B0(n3753), .B1(N153), .C0(
        n3754), .C1(proc_wdata[2]), .Y(n3695) );
  AOI222X4 U274 ( .A0(mem_rdata[33]), .A1(n395), .B0(n3753), .B1(N154), .C0(
        n3754), .C1(proc_wdata[1]), .Y(n3696) );
  AOI222X4 U275 ( .A0(mem_rdata[32]), .A1(n393), .B0(n3753), .B1(N155), .C0(
        n3754), .C1(proc_wdata[0]), .Y(n3697) );
  AOI222X4 U276 ( .A0(mem_rdata[31]), .A1(n395), .B0(n3756), .B1(N156), .C0(
        n3757), .C1(proc_wdata[31]), .Y(n3698) );
  AOI222X4 U277 ( .A0(mem_rdata[30]), .A1(n395), .B0(n3756), .B1(N157), .C0(
        n3757), .C1(proc_wdata[30]), .Y(n3699) );
  AOI222X4 U278 ( .A0(mem_rdata[29]), .A1(n393), .B0(n3756), .B1(N158), .C0(
        n3757), .C1(proc_wdata[29]), .Y(n3700) );
  AOI222X4 U279 ( .A0(mem_rdata[28]), .A1(n395), .B0(n3756), .B1(N159), .C0(
        n3757), .C1(proc_wdata[28]), .Y(n3701) );
  AOI222X4 U280 ( .A0(mem_rdata[27]), .A1(n395), .B0(n3756), .B1(N160), .C0(
        n3757), .C1(proc_wdata[27]), .Y(n3702) );
  AOI222X4 U281 ( .A0(mem_rdata[26]), .A1(n393), .B0(n3756), .B1(N161), .C0(
        n3757), .C1(proc_wdata[26]), .Y(n3703) );
  AOI222X4 U282 ( .A0(mem_rdata[25]), .A1(n396), .B0(n3756), .B1(N162), .C0(
        n3757), .C1(proc_wdata[25]), .Y(n3704) );
  AOI222X4 U283 ( .A0(mem_rdata[24]), .A1(n396), .B0(n3756), .B1(N163), .C0(
        n3757), .C1(proc_wdata[24]), .Y(n3705) );
  AOI222X4 U284 ( .A0(mem_rdata[23]), .A1(n394), .B0(n3756), .B1(N164), .C0(
        n3757), .C1(proc_wdata[23]), .Y(n3706) );
  AOI222X4 U285 ( .A0(mem_rdata[22]), .A1(n396), .B0(n3756), .B1(N165), .C0(
        n3757), .C1(proc_wdata[22]), .Y(n3707) );
  AOI222X4 U286 ( .A0(mem_rdata[21]), .A1(n396), .B0(n3756), .B1(N166), .C0(
        n3757), .C1(proc_wdata[21]), .Y(n3708) );
  AOI222X4 U287 ( .A0(mem_rdata[20]), .A1(n393), .B0(n3756), .B1(N167), .C0(
        n3757), .C1(proc_wdata[20]), .Y(n3709) );
  AOI222X4 U288 ( .A0(mem_rdata[19]), .A1(n396), .B0(n3756), .B1(N168), .C0(
        n3757), .C1(proc_wdata[19]), .Y(n3710) );
  AOI222X4 U289 ( .A0(mem_rdata[18]), .A1(n395), .B0(n3756), .B1(N169), .C0(
        n3757), .C1(proc_wdata[18]), .Y(n3711) );
  AOI222X4 U290 ( .A0(mem_rdata[17]), .A1(n394), .B0(n3756), .B1(N170), .C0(
        n3757), .C1(proc_wdata[17]), .Y(n3712) );
  AOI222X4 U291 ( .A0(mem_rdata[16]), .A1(n396), .B0(n3756), .B1(N171), .C0(
        n3757), .C1(proc_wdata[16]), .Y(n3713) );
  AOI222X4 U292 ( .A0(mem_rdata[15]), .A1(n396), .B0(n3756), .B1(N172), .C0(
        n3757), .C1(proc_wdata[15]), .Y(n3714) );
  AOI222X4 U293 ( .A0(mem_rdata[14]), .A1(n394), .B0(n3756), .B1(N173), .C0(
        n3757), .C1(proc_wdata[14]), .Y(n3715) );
  AOI222X4 U294 ( .A0(mem_rdata[13]), .A1(n396), .B0(n3756), .B1(N174), .C0(
        n3757), .C1(proc_wdata[13]), .Y(n3716) );
  AOI222X4 U295 ( .A0(mem_rdata[12]), .A1(n396), .B0(n3756), .B1(N175), .C0(
        n3757), .C1(proc_wdata[12]), .Y(n3717) );
  AOI222X4 U296 ( .A0(mem_rdata[11]), .A1(n394), .B0(n3756), .B1(N176), .C0(
        n3757), .C1(proc_wdata[11]), .Y(n3718) );
  AOI222X4 U297 ( .A0(mem_rdata[10]), .A1(n395), .B0(n3756), .B1(N177), .C0(
        n3757), .C1(proc_wdata[10]), .Y(n3719) );
  AOI222X4 U298 ( .A0(mem_rdata[9]), .A1(n396), .B0(n3756), .B1(N178), .C0(
        n3757), .C1(proc_wdata[9]), .Y(n3720) );
  AOI222X4 U299 ( .A0(mem_rdata[8]), .A1(n395), .B0(n3756), .B1(N179), .C0(
        n3757), .C1(proc_wdata[8]), .Y(n3721) );
  AOI222X4 U300 ( .A0(mem_rdata[7]), .A1(n396), .B0(n3756), .B1(N180), .C0(
        n3757), .C1(proc_wdata[7]), .Y(n3722) );
  AOI222X4 U301 ( .A0(mem_rdata[6]), .A1(n396), .B0(n3756), .B1(N181), .C0(
        n3757), .C1(proc_wdata[6]), .Y(n3723) );
  AOI222X4 U302 ( .A0(mem_rdata[5]), .A1(n395), .B0(n3756), .B1(N182), .C0(
        n3757), .C1(proc_wdata[5]), .Y(n3724) );
  AOI222X4 U303 ( .A0(mem_rdata[4]), .A1(n396), .B0(n3756), .B1(N183), .C0(
        n3757), .C1(proc_wdata[4]), .Y(n3725) );
  AOI222X4 U304 ( .A0(mem_rdata[3]), .A1(n396), .B0(n3756), .B1(N184), .C0(
        n3757), .C1(proc_wdata[3]), .Y(n3726) );
  AOI222X4 U305 ( .A0(mem_rdata[2]), .A1(n395), .B0(n3756), .B1(N185), .C0(
        n3757), .C1(proc_wdata[2]), .Y(n3727) );
  AOI222X4 U306 ( .A0(mem_rdata[1]), .A1(n396), .B0(n3756), .B1(N186), .C0(
        n3757), .C1(proc_wdata[1]), .Y(n3728) );
  AOI222X4 U307 ( .A0(mem_rdata[0]), .A1(n397), .B0(n3756), .B1(N187), .C0(
        n3757), .C1(proc_wdata[0]), .Y(n3729) );
  INVX12 U308 ( .A(n138), .Y(mem_addr[9]) );
  INVX12 U309 ( .A(n137), .Y(mem_addr[8]) );
  INVX12 U310 ( .A(n136), .Y(mem_addr[7]) );
  INVX12 U311 ( .A(n135), .Y(mem_addr[6]) );
  INVX12 U312 ( .A(n134), .Y(mem_addr[5]) );
  INVX12 U313 ( .A(n133), .Y(mem_addr[4]) );
  INVX12 U314 ( .A(n132), .Y(mem_addr[3]) );
  INVX12 U315 ( .A(n156), .Y(mem_addr[27]) );
  INVX12 U316 ( .A(n155), .Y(mem_addr[26]) );
  INVX12 U317 ( .A(n154), .Y(mem_addr[25]) );
  INVX12 U318 ( .A(n153), .Y(mem_addr[24]) );
  INVX12 U319 ( .A(n152), .Y(mem_addr[23]) );
  INVX12 U320 ( .A(n151), .Y(mem_addr[22]) );
  INVX12 U321 ( .A(n150), .Y(mem_addr[21]) );
  INVX12 U322 ( .A(n149), .Y(mem_addr[20]) );
  INVX12 U323 ( .A(n148), .Y(mem_addr[19]) );
  INVX12 U324 ( .A(n147), .Y(mem_addr[18]) );
  INVX12 U325 ( .A(n146), .Y(mem_addr[17]) );
  INVX12 U326 ( .A(n145), .Y(mem_addr[16]) );
  INVX12 U327 ( .A(n144), .Y(mem_addr[15]) );
  INVX12 U328 ( .A(n143), .Y(mem_addr[14]) );
  INVX12 U329 ( .A(n142), .Y(mem_addr[13]) );
  INVX12 U330 ( .A(n141), .Y(mem_addr[12]) );
  INVX12 U331 ( .A(n140), .Y(mem_addr[11]) );
  INVX12 U332 ( .A(n139), .Y(mem_addr[10]) );
  INVX12 U333 ( .A(n11), .Y(mem_wdata[9]) );
  INVX12 U334 ( .A(n101), .Y(mem_wdata[99]) );
  INVX12 U335 ( .A(n100), .Y(mem_wdata[98]) );
  INVX12 U336 ( .A(n99), .Y(mem_wdata[97]) );
  INVX12 U337 ( .A(n98), .Y(mem_wdata[96]) );
  INVX12 U338 ( .A(n97), .Y(mem_wdata[95]) );
  INVX12 U339 ( .A(n96), .Y(mem_wdata[94]) );
  INVX12 U340 ( .A(n95), .Y(mem_wdata[93]) );
  INVX12 U341 ( .A(n94), .Y(mem_wdata[92]) );
  INVX12 U342 ( .A(n93), .Y(mem_wdata[91]) );
  INVX12 U343 ( .A(n92), .Y(mem_wdata[90]) );
  INVX12 U344 ( .A(n10), .Y(mem_wdata[8]) );
  INVX12 U345 ( .A(n91), .Y(mem_wdata[89]) );
  INVX12 U346 ( .A(n90), .Y(mem_wdata[88]) );
  INVX12 U347 ( .A(n89), .Y(mem_wdata[87]) );
  INVX12 U348 ( .A(n88), .Y(mem_wdata[86]) );
  INVX12 U349 ( .A(n87), .Y(mem_wdata[85]) );
  INVX12 U350 ( .A(n86), .Y(mem_wdata[84]) );
  INVX12 U351 ( .A(n85), .Y(mem_wdata[83]) );
  INVX12 U352 ( .A(n84), .Y(mem_wdata[82]) );
  INVX12 U353 ( .A(n83), .Y(mem_wdata[81]) );
  INVX12 U354 ( .A(n82), .Y(mem_wdata[80]) );
  INVX12 U355 ( .A(n9), .Y(mem_wdata[7]) );
  INVX12 U356 ( .A(n81), .Y(mem_wdata[79]) );
  INVX12 U357 ( .A(n80), .Y(mem_wdata[78]) );
  INVX12 U358 ( .A(n79), .Y(mem_wdata[77]) );
  INVX12 U359 ( .A(n78), .Y(mem_wdata[76]) );
  INVX12 U360 ( .A(n77), .Y(mem_wdata[75]) );
  INVX12 U361 ( .A(n76), .Y(mem_wdata[74]) );
  INVX12 U362 ( .A(n75), .Y(mem_wdata[73]) );
  INVX12 U363 ( .A(n74), .Y(mem_wdata[72]) );
  INVX12 U364 ( .A(n73), .Y(mem_wdata[71]) );
  INVX12 U365 ( .A(n72), .Y(mem_wdata[70]) );
  INVX12 U366 ( .A(n8), .Y(mem_wdata[6]) );
  INVX12 U367 ( .A(n71), .Y(mem_wdata[69]) );
  INVX12 U368 ( .A(n70), .Y(mem_wdata[68]) );
  INVX12 U369 ( .A(n69), .Y(mem_wdata[67]) );
  INVX12 U370 ( .A(n68), .Y(mem_wdata[66]) );
  INVX12 U371 ( .A(n67), .Y(mem_wdata[65]) );
  INVX12 U372 ( .A(n66), .Y(mem_wdata[64]) );
  INVX12 U373 ( .A(n65), .Y(mem_wdata[63]) );
  INVX12 U374 ( .A(n64), .Y(mem_wdata[62]) );
  INVX12 U375 ( .A(n63), .Y(mem_wdata[61]) );
  INVX12 U376 ( .A(n62), .Y(mem_wdata[60]) );
  INVX12 U377 ( .A(n7), .Y(mem_wdata[5]) );
  INVX12 U378 ( .A(n61), .Y(mem_wdata[59]) );
  INVX12 U379 ( .A(n60), .Y(mem_wdata[58]) );
  INVX12 U380 ( .A(n59), .Y(mem_wdata[57]) );
  INVX12 U381 ( .A(n58), .Y(mem_wdata[56]) );
  INVX12 U382 ( .A(n57), .Y(mem_wdata[55]) );
  INVX12 U383 ( .A(n56), .Y(mem_wdata[54]) );
  INVX12 U384 ( .A(n55), .Y(mem_wdata[53]) );
  INVX12 U385 ( .A(n54), .Y(mem_wdata[52]) );
  INVX12 U386 ( .A(n53), .Y(mem_wdata[51]) );
  INVX12 U387 ( .A(n52), .Y(mem_wdata[50]) );
  INVX12 U388 ( .A(n6), .Y(mem_wdata[4]) );
  INVX12 U389 ( .A(n51), .Y(mem_wdata[49]) );
  INVX12 U390 ( .A(n50), .Y(mem_wdata[48]) );
  INVX12 U391 ( .A(n49), .Y(mem_wdata[47]) );
  INVX12 U392 ( .A(n48), .Y(mem_wdata[46]) );
  INVX12 U393 ( .A(n47), .Y(mem_wdata[45]) );
  INVX12 U394 ( .A(n46), .Y(mem_wdata[44]) );
  INVX12 U395 ( .A(n45), .Y(mem_wdata[43]) );
  INVX12 U396 ( .A(n44), .Y(mem_wdata[42]) );
  INVX12 U397 ( .A(n43), .Y(mem_wdata[41]) );
  INVX12 U398 ( .A(n42), .Y(mem_wdata[40]) );
  INVX12 U399 ( .A(n5), .Y(mem_wdata[3]) );
  INVX12 U400 ( .A(n41), .Y(mem_wdata[39]) );
  INVX12 U401 ( .A(n40), .Y(mem_wdata[38]) );
  INVX12 U402 ( .A(n39), .Y(mem_wdata[37]) );
  INVX12 U403 ( .A(n38), .Y(mem_wdata[36]) );
  INVX12 U404 ( .A(n37), .Y(mem_wdata[35]) );
  INVX12 U405 ( .A(n36), .Y(mem_wdata[34]) );
  INVX12 U406 ( .A(n35), .Y(mem_wdata[33]) );
  INVX12 U407 ( .A(n34), .Y(mem_wdata[32]) );
  INVX12 U408 ( .A(n33), .Y(mem_wdata[31]) );
  INVX12 U409 ( .A(n32), .Y(mem_wdata[30]) );
  INVX12 U410 ( .A(n4), .Y(mem_wdata[2]) );
  INVX12 U411 ( .A(n31), .Y(mem_wdata[29]) );
  INVX12 U412 ( .A(n30), .Y(mem_wdata[28]) );
  INVX12 U413 ( .A(n29), .Y(mem_wdata[27]) );
  INVX12 U414 ( .A(n28), .Y(mem_wdata[26]) );
  INVX12 U415 ( .A(n27), .Y(mem_wdata[25]) );
  INVX12 U416 ( .A(n26), .Y(mem_wdata[24]) );
  INVX12 U417 ( .A(n25), .Y(mem_wdata[23]) );
  INVX12 U418 ( .A(n24), .Y(mem_wdata[22]) );
  INVX12 U419 ( .A(n23), .Y(mem_wdata[21]) );
  INVX12 U420 ( .A(n22), .Y(mem_wdata[20]) );
  INVX12 U421 ( .A(n3), .Y(mem_wdata[1]) );
  INVX12 U422 ( .A(n21), .Y(mem_wdata[19]) );
  INVX12 U423 ( .A(n20), .Y(mem_wdata[18]) );
  INVX12 U424 ( .A(n19), .Y(mem_wdata[17]) );
  INVX12 U425 ( .A(n18), .Y(mem_wdata[16]) );
  INVX12 U426 ( .A(n17), .Y(mem_wdata[15]) );
  INVX12 U427 ( .A(n16), .Y(mem_wdata[14]) );
  INVX12 U428 ( .A(n15), .Y(mem_wdata[13]) );
  INVX12 U429 ( .A(n14), .Y(mem_wdata[12]) );
  INVX12 U430 ( .A(n129), .Y(mem_wdata[127]) );
  INVX12 U431 ( .A(n128), .Y(mem_wdata[126]) );
  INVX12 U432 ( .A(n127), .Y(mem_wdata[125]) );
  INVX12 U433 ( .A(n126), .Y(mem_wdata[124]) );
  INVX12 U434 ( .A(n125), .Y(mem_wdata[123]) );
  INVX12 U435 ( .A(n124), .Y(mem_wdata[122]) );
  INVX12 U436 ( .A(n123), .Y(mem_wdata[121]) );
  INVX12 U437 ( .A(n122), .Y(mem_wdata[120]) );
  INVX12 U438 ( .A(n13), .Y(mem_wdata[11]) );
  INVX12 U439 ( .A(n121), .Y(mem_wdata[119]) );
  INVX12 U440 ( .A(n120), .Y(mem_wdata[118]) );
  INVX12 U441 ( .A(n119), .Y(mem_wdata[117]) );
  INVX12 U442 ( .A(n118), .Y(mem_wdata[116]) );
  INVX12 U443 ( .A(n117), .Y(mem_wdata[115]) );
  INVX12 U444 ( .A(n116), .Y(mem_wdata[114]) );
  INVX12 U445 ( .A(n115), .Y(mem_wdata[113]) );
  INVX12 U446 ( .A(n114), .Y(mem_wdata[112]) );
  INVX12 U447 ( .A(n113), .Y(mem_wdata[111]) );
  INVX12 U448 ( .A(n112), .Y(mem_wdata[110]) );
  INVX12 U449 ( .A(n12), .Y(mem_wdata[10]) );
  INVX12 U450 ( .A(n111), .Y(mem_wdata[109]) );
  INVX12 U451 ( .A(n110), .Y(mem_wdata[108]) );
  INVX12 U452 ( .A(n109), .Y(mem_wdata[107]) );
  INVX12 U453 ( .A(n108), .Y(mem_wdata[106]) );
  INVX12 U454 ( .A(n107), .Y(mem_wdata[105]) );
  INVX12 U455 ( .A(n106), .Y(mem_wdata[104]) );
  INVX12 U456 ( .A(n105), .Y(mem_wdata[103]) );
  INVX12 U457 ( .A(n104), .Y(mem_wdata[102]) );
  INVX12 U458 ( .A(n103), .Y(mem_wdata[101]) );
  INVX12 U459 ( .A(n102), .Y(mem_wdata[100]) );
  INVX12 U460 ( .A(n2), .Y(mem_wdata[0]) );
  INVX12 U461 ( .A(n1), .Y(mem_addr[2]) );
  INVX12 U462 ( .A(n131), .Y(mem_addr[1]) );
  INVX12 U463 ( .A(n130), .Y(mem_addr[0]) );
  CLKINVX1 U464 ( .A(n6281), .Y(n313) );
  INVX16 U465 ( .A(n313), .Y(mem_read) );
  CLKINVX2 U466 ( .A(proc_addr[1]), .Y(n3573) );
  NAND3X6 U467 ( .A(n3572), .B(n3573), .C(n3571), .Y(n3412) );
  NOR3X6 U468 ( .A(n3573), .B(n3572), .C(n3739), .Y(n3746) );
  CLKINVX2 U469 ( .A(proc_addr[0]), .Y(n3572) );
  AOI211X1 U470 ( .A0(n3762), .A1(N34), .B0(n3571), .C0(n3404), .Y(n3744) );
  INVX6 U471 ( .A(n3752), .Y(n3751) );
  INVX6 U472 ( .A(n3758), .Y(n3756) );
  INVX6 U473 ( .A(n3755), .Y(n3753) );
  NAND3X6 U474 ( .A(proc_addr[0]), .B(n3571), .C(proc_addr[1]), .Y(n3414) );
  AOI22X2 U475 ( .A0(proc_addr[5]), .A1(n398), .B0(n3742), .B1(N59), .Y(n3601)
         );
  AOI22X2 U476 ( .A0(proc_addr[6]), .A1(n392), .B0(n3742), .B1(N58), .Y(n3600)
         );
  AOI22X2 U477 ( .A0(proc_addr[7]), .A1(n392), .B0(n3742), .B1(N57), .Y(n3599)
         );
  AOI22X2 U478 ( .A0(proc_addr[8]), .A1(n392), .B0(n3742), .B1(N56), .Y(n3598)
         );
  AOI22X2 U479 ( .A0(proc_addr[9]), .A1(n392), .B0(n3742), .B1(N55), .Y(n3597)
         );
  AOI22X2 U480 ( .A0(proc_addr[10]), .A1(n392), .B0(n3742), .B1(N54), .Y(n3596) );
  NAND3X6 U481 ( .A(n3743), .B(n3739), .C(n3744), .Y(n3742) );
  NAND3X6 U482 ( .A(n3571), .B(n3572), .C(proc_addr[1]), .Y(n3407) );
  NAND3X6 U483 ( .A(n3571), .B(n3573), .C(proc_addr[0]), .Y(n3409) );
  NOR2X2 U484 ( .A(n3763), .B(n3760), .Y(n3571) );
  INVX6 U485 ( .A(n3747), .Y(n3745) );
  NOR3X6 U486 ( .A(proc_addr[0]), .B(proc_addr[1]), .C(n3739), .Y(n3757) );
  OAI221X1 U487 ( .A0(n3406), .A1(n3743), .B0(mem_ready), .B1(n3761), .C0(
        n3744), .Y(n3748) );
  AOI211X4 U488 ( .A0(proc_read), .A1(mem_ready), .B0(n3737), .C0(N33), .Y(
        n3574) );
  NOR3X6 U489 ( .A(n3572), .B(proc_addr[1]), .C(n3739), .Y(n3754) );
  NOR3X6 U490 ( .A(n3573), .B(proc_addr[0]), .C(n3739), .Y(n3750) );
  INVX3 U491 ( .A(n3737), .Y(n3739) );
  OA22XL U492 ( .A0(n3412), .A1(n3539), .B0(n3414), .B1(n3540), .Y(n3538) );
  OA22XL U493 ( .A0(n3412), .A1(n3524), .B0(n3414), .B1(n3525), .Y(n3523) );
  OA22XL U494 ( .A0(n3412), .A1(n3519), .B0(n3414), .B1(n3520), .Y(n3518) );
  OA22XL U495 ( .A0(n3412), .A1(n3509), .B0(n3414), .B1(n3510), .Y(n3508) );
  OA22XL U496 ( .A0(n3412), .A1(n3494), .B0(n3414), .B1(n3495), .Y(n3493) );
  OA22XL U497 ( .A0(n3412), .A1(n3489), .B0(n3414), .B1(n3490), .Y(n3488) );
  OA22XL U498 ( .A0(n3412), .A1(n3484), .B0(n3414), .B1(n3485), .Y(n3483) );
  OA22XL U499 ( .A0(n3412), .A1(n3464), .B0(n3414), .B1(n3465), .Y(n3463) );
  OA22XL U500 ( .A0(n3412), .A1(n3569), .B0(n3414), .B1(n3570), .Y(n3568) );
  OA22XL U501 ( .A0(n3412), .A1(n3514), .B0(n3414), .B1(n3515), .Y(n3513) );
  OA22XL U502 ( .A0(n3412), .A1(n3459), .B0(n3414), .B1(n3460), .Y(n3458) );
  OA22XL U503 ( .A0(n3412), .A1(n3444), .B0(n3414), .B1(n3445), .Y(n3443) );
  OA22XL U504 ( .A0(n3412), .A1(n3439), .B0(n3414), .B1(n3440), .Y(n3438) );
  OA22XL U505 ( .A0(n3412), .A1(n3434), .B0(n3414), .B1(n3435), .Y(n3433) );
  OA22XL U506 ( .A0(n3412), .A1(n3429), .B0(n3414), .B1(n3430), .Y(n3428) );
  OA22XL U507 ( .A0(n3412), .A1(n3424), .B0(n3414), .B1(n3425), .Y(n3423) );
  OA22XL U508 ( .A0(n3412), .A1(n3419), .B0(n3414), .B1(n3420), .Y(n3418) );
  OA22XL U509 ( .A0(n3412), .A1(n3413), .B0(n3414), .B1(n3415), .Y(n3411) );
  OA22XL U510 ( .A0(n3412), .A1(n3564), .B0(n3414), .B1(n3565), .Y(n3563) );
  OA22XL U511 ( .A0(n3412), .A1(n3559), .B0(n3414), .B1(n3560), .Y(n3558) );
  OA22XL U512 ( .A0(n3412), .A1(n3554), .B0(n3414), .B1(n3555), .Y(n3553) );
  OA22XL U513 ( .A0(n3412), .A1(n3549), .B0(n3414), .B1(n3550), .Y(n3548) );
  OA22XL U514 ( .A0(n3412), .A1(n3544), .B0(n3414), .B1(n3545), .Y(n3543) );
  OA22XL U515 ( .A0(n3412), .A1(n3534), .B0(n3414), .B1(n3535), .Y(n3533) );
  OA22XL U516 ( .A0(n3412), .A1(n3529), .B0(n3414), .B1(n3530), .Y(n3528) );
  OA22XL U517 ( .A0(n3412), .A1(n3504), .B0(n3414), .B1(n3505), .Y(n3503) );
  OA22XL U518 ( .A0(n3412), .A1(n3499), .B0(n3414), .B1(n3500), .Y(n3498) );
  OA22XL U519 ( .A0(n3412), .A1(n3479), .B0(n3414), .B1(n3480), .Y(n3478) );
  OA22XL U520 ( .A0(n3412), .A1(n3474), .B0(n3414), .B1(n3475), .Y(n3473) );
  OA22XL U521 ( .A0(n3412), .A1(n3469), .B0(n3414), .B1(n3470), .Y(n3468) );
  OA22XL U522 ( .A0(n3412), .A1(n3454), .B0(n3414), .B1(n3455), .Y(n3453) );
  OA22XL U523 ( .A0(n3412), .A1(n3449), .B0(n3414), .B1(n3450), .Y(n3448) );
  AND2X2 U524 ( .A(n3738), .B(n3739), .Y(n3576) );
  MXI2XL U525 ( .A(n6280), .B(n3729), .S0(n382), .Y(n5040) );
  MXI2XL U526 ( .A(n6279), .B(n3728), .S0(n382), .Y(n5039) );
  MXI2XL U527 ( .A(n6278), .B(n3727), .S0(n382), .Y(n5038) );
  MXI2XL U528 ( .A(n6277), .B(n3726), .S0(n382), .Y(n5037) );
  MXI2XL U529 ( .A(n6276), .B(n3725), .S0(n382), .Y(n5036) );
  MXI2XL U530 ( .A(n6275), .B(n3724), .S0(n382), .Y(n5035) );
  MXI2XL U531 ( .A(n6274), .B(n3723), .S0(n382), .Y(n5034) );
  MXI2XL U532 ( .A(n6273), .B(n3722), .S0(n382), .Y(n5033) );
  MXI2XL U533 ( .A(n6272), .B(n3721), .S0(n382), .Y(n5032) );
  MXI2XL U534 ( .A(n6271), .B(n3720), .S0(n382), .Y(n5031) );
  MXI2XL U535 ( .A(n6270), .B(n3719), .S0(n382), .Y(n5030) );
  MXI2XL U536 ( .A(n6269), .B(n3718), .S0(n382), .Y(n5029) );
  MXI2XL U537 ( .A(n6268), .B(n3717), .S0(n382), .Y(n5028) );
  MXI2XL U538 ( .A(n6267), .B(n3716), .S0(n383), .Y(n5027) );
  MXI2XL U539 ( .A(n6266), .B(n3715), .S0(n383), .Y(n5026) );
  MXI2XL U540 ( .A(n6265), .B(n3714), .S0(n383), .Y(n5025) );
  MXI2XL U541 ( .A(n6264), .B(n3713), .S0(n383), .Y(n5024) );
  MXI2XL U542 ( .A(n6263), .B(n3712), .S0(n383), .Y(n5023) );
  MXI2XL U543 ( .A(n6262), .B(n3711), .S0(n383), .Y(n5022) );
  MXI2XL U544 ( .A(n6261), .B(n3710), .S0(n383), .Y(n5021) );
  MXI2XL U545 ( .A(n6260), .B(n3709), .S0(n383), .Y(n5020) );
  MXI2XL U546 ( .A(n6259), .B(n3708), .S0(n383), .Y(n5019) );
  MXI2XL U547 ( .A(n6258), .B(n3707), .S0(n383), .Y(n5018) );
  MXI2XL U548 ( .A(n6257), .B(n3706), .S0(n383), .Y(n5017) );
  MXI2XL U549 ( .A(n6256), .B(n3705), .S0(n383), .Y(n5016) );
  MXI2XL U550 ( .A(n6255), .B(n3704), .S0(n383), .Y(n5015) );
  MXI2XL U551 ( .A(n6254), .B(n3703), .S0(n384), .Y(n5014) );
  MXI2XL U552 ( .A(n6253), .B(n3702), .S0(n384), .Y(n5013) );
  MXI2XL U553 ( .A(n6252), .B(n3701), .S0(n384), .Y(n5012) );
  MXI2XL U554 ( .A(n6251), .B(n3700), .S0(n384), .Y(n5011) );
  MXI2XL U555 ( .A(n6250), .B(n3699), .S0(n384), .Y(n5010) );
  MXI2XL U556 ( .A(n6249), .B(n3698), .S0(n384), .Y(n5009) );
  MXI2XL U557 ( .A(n6248), .B(n3697), .S0(n384), .Y(n5008) );
  MXI2XL U558 ( .A(n6247), .B(n3696), .S0(n384), .Y(n5007) );
  MXI2XL U559 ( .A(n6246), .B(n3695), .S0(n384), .Y(n5006) );
  MXI2XL U560 ( .A(n6245), .B(n3694), .S0(n384), .Y(n5005) );
  MXI2XL U561 ( .A(n6244), .B(n3693), .S0(n384), .Y(n5004) );
  MXI2XL U562 ( .A(n6243), .B(n3692), .S0(n384), .Y(n5003) );
  MXI2XL U563 ( .A(n6242), .B(n3691), .S0(n384), .Y(n5002) );
  MXI2XL U564 ( .A(n6241), .B(n3690), .S0(n385), .Y(n5001) );
  MXI2XL U565 ( .A(n6240), .B(n3689), .S0(n385), .Y(n5000) );
  MXI2XL U566 ( .A(n6239), .B(n3688), .S0(n385), .Y(n4999) );
  MXI2XL U567 ( .A(n6238), .B(n3687), .S0(n385), .Y(n4998) );
  MXI2XL U568 ( .A(n6237), .B(n3686), .S0(n385), .Y(n4997) );
  MXI2XL U569 ( .A(n6236), .B(n3685), .S0(n385), .Y(n4996) );
  MXI2XL U570 ( .A(n6235), .B(n3684), .S0(n385), .Y(n4995) );
  MXI2XL U571 ( .A(n6234), .B(n3683), .S0(n385), .Y(n4994) );
  MXI2XL U572 ( .A(n6233), .B(n3682), .S0(n385), .Y(n4993) );
  MXI2XL U573 ( .A(n6232), .B(n3681), .S0(n385), .Y(n4992) );
  MXI2XL U574 ( .A(n6231), .B(n3680), .S0(n385), .Y(n4991) );
  MXI2XL U575 ( .A(n6230), .B(n3679), .S0(n385), .Y(n4990) );
  MXI2XL U576 ( .A(n6229), .B(n3678), .S0(n385), .Y(n4989) );
  MXI2XL U577 ( .A(n6228), .B(n3677), .S0(n386), .Y(n4988) );
  MXI2XL U578 ( .A(n6227), .B(n3676), .S0(n386), .Y(n4987) );
  MXI2XL U579 ( .A(n6226), .B(n3675), .S0(n386), .Y(n4986) );
  MXI2XL U580 ( .A(n6225), .B(n3674), .S0(n386), .Y(n4985) );
  MXI2XL U581 ( .A(n6224), .B(n3673), .S0(n386), .Y(n4984) );
  MXI2XL U582 ( .A(n6223), .B(n3672), .S0(n386), .Y(n4983) );
  MXI2XL U583 ( .A(n6222), .B(n3671), .S0(n386), .Y(n4982) );
  MXI2XL U584 ( .A(n6221), .B(n3670), .S0(n386), .Y(n4981) );
  MXI2XL U585 ( .A(n6220), .B(n3669), .S0(n386), .Y(n4980) );
  MXI2XL U586 ( .A(n6219), .B(n3668), .S0(n386), .Y(n4979) );
  MXI2XL U587 ( .A(n6218), .B(n3667), .S0(n386), .Y(n4978) );
  MXI2XL U588 ( .A(n6217), .B(n3666), .S0(n386), .Y(n4977) );
  MXI2XL U589 ( .A(n6184), .B(n3633), .S0(n3736), .Y(n4944) );
  MXI2XL U590 ( .A(n6183), .B(n3632), .S0(n384), .Y(n4943) );
  MXI2XL U591 ( .A(n6182), .B(n3631), .S0(n388), .Y(n4942) );
  MXI2XL U592 ( .A(n6181), .B(n3630), .S0(n385), .Y(n4941) );
  MXI2XL U593 ( .A(n6180), .B(n3629), .S0(n389), .Y(n4940) );
  MXI2XL U594 ( .A(n6179), .B(n3628), .S0(n382), .Y(n4939) );
  MXI2XL U595 ( .A(n6178), .B(n3627), .S0(n383), .Y(n4938) );
  MXI2XL U596 ( .A(n6177), .B(n3626), .S0(n386), .Y(n4937) );
  MXI2XL U597 ( .A(n6176), .B(n3625), .S0(n389), .Y(n4936) );
  MXI2XL U598 ( .A(n6175), .B(n3624), .S0(n389), .Y(n4935) );
  MXI2XL U599 ( .A(n6174), .B(n3623), .S0(n389), .Y(n4934) );
  MXI2XL U600 ( .A(n6173), .B(n3622), .S0(n389), .Y(n4933) );
  MXI2XL U601 ( .A(n6172), .B(n3621), .S0(n389), .Y(n4932) );
  MXI2XL U602 ( .A(n6171), .B(n3620), .S0(n389), .Y(n4931) );
  MXI2XL U603 ( .A(n6170), .B(n3619), .S0(n389), .Y(n4930) );
  MXI2XL U604 ( .A(n6169), .B(n3618), .S0(n389), .Y(n4929) );
  MXI2XL U605 ( .A(n6168), .B(n3617), .S0(n389), .Y(n4928) );
  MXI2XL U606 ( .A(n6167), .B(n3616), .S0(n389), .Y(n4927) );
  MXI2XL U607 ( .A(n6166), .B(n3615), .S0(n389), .Y(n4926) );
  MXI2XL U608 ( .A(n6165), .B(n3614), .S0(n389), .Y(n4925) );
  MXI2XL U609 ( .A(n6164), .B(n3613), .S0(n389), .Y(n4924) );
  MXI2XL U610 ( .A(n6163), .B(n3612), .S0(n383), .Y(n4923) );
  MXI2XL U611 ( .A(n6162), .B(n3611), .S0(n386), .Y(n4922) );
  MXI2XL U612 ( .A(n6161), .B(n3610), .S0(n390), .Y(n4921) );
  MXI2XL U613 ( .A(n6160), .B(n3609), .S0(n3736), .Y(n4920) );
  MXI2XL U614 ( .A(n6159), .B(n3608), .S0(n387), .Y(n4919) );
  MXI2XL U615 ( .A(n6158), .B(n3607), .S0(n384), .Y(n4918) );
  MXI2XL U616 ( .A(n6157), .B(n3606), .S0(n388), .Y(n4917) );
  MXI2XL U617 ( .A(n6156), .B(n3605), .S0(n385), .Y(n4916) );
  MXI2XL U618 ( .A(n6155), .B(n3604), .S0(n389), .Y(n4915) );
  MXI2XL U619 ( .A(n6154), .B(n3603), .S0(n382), .Y(n4914) );
  MXI2XL U620 ( .A(n6153), .B(n3602), .S0(n383), .Y(n4913) );
  MXI2XL U621 ( .A(n6125), .B(n3729), .S0(n373), .Y(n4885) );
  MXI2XL U622 ( .A(n6124), .B(n3728), .S0(n373), .Y(n4884) );
  MXI2XL U623 ( .A(n6123), .B(n3727), .S0(n373), .Y(n4883) );
  MXI2XL U624 ( .A(n6122), .B(n3726), .S0(n373), .Y(n4882) );
  MXI2XL U625 ( .A(n6121), .B(n3725), .S0(n373), .Y(n4881) );
  MXI2XL U626 ( .A(n6120), .B(n3724), .S0(n373), .Y(n4880) );
  MXI2XL U627 ( .A(n6119), .B(n3723), .S0(n373), .Y(n4879) );
  MXI2XL U628 ( .A(n6118), .B(n3722), .S0(n373), .Y(n4878) );
  MXI2XL U629 ( .A(n6117), .B(n3721), .S0(n373), .Y(n4877) );
  MXI2XL U630 ( .A(n6116), .B(n3720), .S0(n373), .Y(n4876) );
  MXI2XL U631 ( .A(n6115), .B(n3719), .S0(n373), .Y(n4875) );
  MXI2XL U632 ( .A(n6114), .B(n3718), .S0(n373), .Y(n4874) );
  MXI2XL U633 ( .A(n6113), .B(n3717), .S0(n373), .Y(n4873) );
  MXI2XL U634 ( .A(n6112), .B(n3716), .S0(n374), .Y(n4872) );
  MXI2XL U635 ( .A(n6111), .B(n3715), .S0(n374), .Y(n4871) );
  MXI2XL U636 ( .A(n6110), .B(n3714), .S0(n374), .Y(n4870) );
  MXI2XL U637 ( .A(n6109), .B(n3713), .S0(n374), .Y(n4869) );
  MXI2XL U638 ( .A(n6108), .B(n3712), .S0(n374), .Y(n4868) );
  MXI2XL U639 ( .A(n6107), .B(n3711), .S0(n374), .Y(n4867) );
  MXI2XL U640 ( .A(n6106), .B(n3710), .S0(n374), .Y(n4866) );
  MXI2XL U641 ( .A(n6105), .B(n3709), .S0(n374), .Y(n4865) );
  MXI2XL U642 ( .A(n6104), .B(n3708), .S0(n374), .Y(n4864) );
  MXI2XL U643 ( .A(n6103), .B(n3707), .S0(n374), .Y(n4863) );
  MXI2XL U644 ( .A(n6102), .B(n3706), .S0(n374), .Y(n4862) );
  MXI2XL U645 ( .A(n6101), .B(n3705), .S0(n374), .Y(n4861) );
  MXI2XL U646 ( .A(n6100), .B(n3704), .S0(n374), .Y(n4860) );
  MXI2XL U647 ( .A(n6099), .B(n3703), .S0(n375), .Y(n4859) );
  MXI2XL U648 ( .A(n6098), .B(n3702), .S0(n375), .Y(n4858) );
  MXI2XL U649 ( .A(n6097), .B(n3701), .S0(n375), .Y(n4857) );
  MXI2XL U650 ( .A(n6096), .B(n3700), .S0(n375), .Y(n4856) );
  MXI2XL U651 ( .A(n6095), .B(n3699), .S0(n375), .Y(n4855) );
  MXI2XL U652 ( .A(n6094), .B(n3698), .S0(n375), .Y(n4854) );
  MXI2XL U653 ( .A(n6093), .B(n3697), .S0(n375), .Y(n4853) );
  MXI2XL U654 ( .A(n6092), .B(n3696), .S0(n375), .Y(n4852) );
  MXI2XL U655 ( .A(n6091), .B(n3695), .S0(n375), .Y(n4851) );
  MXI2XL U656 ( .A(n6090), .B(n3694), .S0(n375), .Y(n4850) );
  MXI2XL U657 ( .A(n6089), .B(n3693), .S0(n375), .Y(n4849) );
  MXI2XL U658 ( .A(n6088), .B(n3692), .S0(n375), .Y(n4848) );
  MXI2XL U659 ( .A(n6087), .B(n3691), .S0(n375), .Y(n4847) );
  MXI2XL U660 ( .A(n6086), .B(n3690), .S0(n376), .Y(n4846) );
  MXI2XL U661 ( .A(n6085), .B(n3689), .S0(n376), .Y(n4845) );
  MXI2XL U662 ( .A(n6084), .B(n3688), .S0(n376), .Y(n4844) );
  MXI2XL U663 ( .A(n6083), .B(n3687), .S0(n376), .Y(n4843) );
  MXI2XL U664 ( .A(n6082), .B(n3686), .S0(n376), .Y(n4842) );
  MXI2XL U665 ( .A(n6081), .B(n3685), .S0(n376), .Y(n4841) );
  MXI2XL U666 ( .A(n6080), .B(n3684), .S0(n376), .Y(n4840) );
  MXI2XL U667 ( .A(n6079), .B(n3683), .S0(n376), .Y(n4839) );
  MXI2XL U668 ( .A(n6078), .B(n3682), .S0(n376), .Y(n4838) );
  MXI2XL U669 ( .A(n6077), .B(n3681), .S0(n376), .Y(n4837) );
  MXI2XL U670 ( .A(n6076), .B(n3680), .S0(n376), .Y(n4836) );
  MXI2XL U671 ( .A(n6075), .B(n3679), .S0(n376), .Y(n4835) );
  MXI2XL U672 ( .A(n6074), .B(n3678), .S0(n376), .Y(n4834) );
  MXI2XL U673 ( .A(n6073), .B(n3677), .S0(n377), .Y(n4833) );
  MXI2XL U674 ( .A(n6072), .B(n3676), .S0(n377), .Y(n4832) );
  MXI2XL U675 ( .A(n6071), .B(n3675), .S0(n377), .Y(n4831) );
  MXI2XL U676 ( .A(n6070), .B(n3674), .S0(n377), .Y(n4830) );
  MXI2XL U677 ( .A(n6069), .B(n3673), .S0(n377), .Y(n4829) );
  MXI2XL U678 ( .A(n6068), .B(n3672), .S0(n377), .Y(n4828) );
  MXI2XL U679 ( .A(n6067), .B(n3671), .S0(n377), .Y(n4827) );
  MXI2XL U680 ( .A(n6066), .B(n3670), .S0(n377), .Y(n4826) );
  MXI2XL U681 ( .A(n6065), .B(n3669), .S0(n377), .Y(n4825) );
  MXI2XL U682 ( .A(n6064), .B(n3668), .S0(n377), .Y(n4824) );
  MXI2XL U683 ( .A(n6063), .B(n3667), .S0(n377), .Y(n4823) );
  MXI2XL U684 ( .A(n6062), .B(n3666), .S0(n377), .Y(n4822) );
  MXI2XL U685 ( .A(n6029), .B(n3633), .S0(n3735), .Y(n4789) );
  MXI2XL U686 ( .A(n6028), .B(n3632), .S0(n375), .Y(n4788) );
  MXI2XL U687 ( .A(n6027), .B(n3631), .S0(n379), .Y(n4787) );
  MXI2XL U688 ( .A(n6026), .B(n3630), .S0(n376), .Y(n4786) );
  MXI2XL U689 ( .A(n6025), .B(n3629), .S0(n380), .Y(n4785) );
  MXI2XL U690 ( .A(n6024), .B(n3628), .S0(n373), .Y(n4784) );
  MXI2XL U691 ( .A(n6023), .B(n3627), .S0(n374), .Y(n4783) );
  MXI2XL U692 ( .A(n6022), .B(n3626), .S0(n377), .Y(n4782) );
  MXI2XL U693 ( .A(n6021), .B(n3625), .S0(n380), .Y(n4781) );
  MXI2XL U694 ( .A(n6020), .B(n3624), .S0(n380), .Y(n4780) );
  MXI2XL U695 ( .A(n6019), .B(n3623), .S0(n380), .Y(n4779) );
  MXI2XL U696 ( .A(n6018), .B(n3622), .S0(n380), .Y(n4778) );
  MXI2XL U697 ( .A(n6017), .B(n3621), .S0(n380), .Y(n4777) );
  MXI2XL U698 ( .A(n6016), .B(n3620), .S0(n380), .Y(n4776) );
  MXI2XL U699 ( .A(n6015), .B(n3619), .S0(n380), .Y(n4775) );
  MXI2XL U700 ( .A(n6014), .B(n3618), .S0(n380), .Y(n4774) );
  MXI2XL U701 ( .A(n6013), .B(n3617), .S0(n380), .Y(n4773) );
  MXI2XL U702 ( .A(n6012), .B(n3616), .S0(n380), .Y(n4772) );
  MXI2XL U703 ( .A(n6011), .B(n3615), .S0(n380), .Y(n4771) );
  MXI2XL U704 ( .A(n6010), .B(n3614), .S0(n380), .Y(n4770) );
  MXI2XL U705 ( .A(n6009), .B(n3613), .S0(n380), .Y(n4769) );
  MXI2XL U706 ( .A(n6008), .B(n3612), .S0(n374), .Y(n4768) );
  MXI2XL U707 ( .A(n6007), .B(n3611), .S0(n377), .Y(n4767) );
  MXI2XL U708 ( .A(n6006), .B(n3610), .S0(n381), .Y(n4766) );
  MXI2XL U709 ( .A(n6005), .B(n3609), .S0(n3735), .Y(n4765) );
  MXI2XL U710 ( .A(n6004), .B(n3608), .S0(n378), .Y(n4764) );
  MXI2XL U711 ( .A(n6003), .B(n3607), .S0(n375), .Y(n4763) );
  MXI2XL U712 ( .A(n6002), .B(n3606), .S0(n379), .Y(n4762) );
  MXI2XL U713 ( .A(n6001), .B(n3605), .S0(n376), .Y(n4761) );
  MXI2XL U714 ( .A(n6000), .B(n3604), .S0(n380), .Y(n4760) );
  MXI2XL U715 ( .A(n5999), .B(n3603), .S0(n373), .Y(n4759) );
  MXI2XL U716 ( .A(n5998), .B(n3602), .S0(n374), .Y(n4758) );
  MXI2XL U717 ( .A(n5970), .B(n3729), .S0(n364), .Y(n4730) );
  MXI2XL U718 ( .A(n5969), .B(n3728), .S0(n364), .Y(n4729) );
  MXI2XL U719 ( .A(n5968), .B(n3727), .S0(n364), .Y(n4728) );
  MXI2XL U720 ( .A(n5967), .B(n3726), .S0(n364), .Y(n4727) );
  MXI2XL U721 ( .A(n5966), .B(n3725), .S0(n364), .Y(n4726) );
  MXI2XL U722 ( .A(n5965), .B(n3724), .S0(n364), .Y(n4725) );
  MXI2XL U723 ( .A(n5964), .B(n3723), .S0(n364), .Y(n4724) );
  MXI2XL U724 ( .A(n5963), .B(n3722), .S0(n364), .Y(n4723) );
  MXI2XL U725 ( .A(n5962), .B(n3721), .S0(n364), .Y(n4722) );
  MXI2XL U726 ( .A(n5961), .B(n3720), .S0(n364), .Y(n4721) );
  MXI2XL U727 ( .A(n5960), .B(n3719), .S0(n364), .Y(n4720) );
  MXI2XL U728 ( .A(n5959), .B(n3718), .S0(n364), .Y(n4719) );
  MXI2XL U729 ( .A(n5958), .B(n3717), .S0(n364), .Y(n4718) );
  MXI2XL U730 ( .A(n5957), .B(n3716), .S0(n365), .Y(n4717) );
  MXI2XL U731 ( .A(n5956), .B(n3715), .S0(n365), .Y(n4716) );
  MXI2XL U732 ( .A(n5955), .B(n3714), .S0(n365), .Y(n4715) );
  MXI2XL U733 ( .A(n5954), .B(n3713), .S0(n365), .Y(n4714) );
  MXI2XL U734 ( .A(n5953), .B(n3712), .S0(n365), .Y(n4713) );
  MXI2XL U735 ( .A(n5952), .B(n3711), .S0(n365), .Y(n4712) );
  MXI2XL U736 ( .A(n5951), .B(n3710), .S0(n365), .Y(n4711) );
  MXI2XL U737 ( .A(n5950), .B(n3709), .S0(n365), .Y(n4710) );
  MXI2XL U738 ( .A(n5949), .B(n3708), .S0(n365), .Y(n4709) );
  MXI2XL U739 ( .A(n5948), .B(n3707), .S0(n365), .Y(n4708) );
  MXI2XL U740 ( .A(n5947), .B(n3706), .S0(n365), .Y(n4707) );
  MXI2XL U741 ( .A(n5946), .B(n3705), .S0(n365), .Y(n4706) );
  MXI2XL U742 ( .A(n5945), .B(n3704), .S0(n365), .Y(n4705) );
  MXI2XL U743 ( .A(n5944), .B(n3703), .S0(n366), .Y(n4704) );
  MXI2XL U744 ( .A(n5943), .B(n3702), .S0(n366), .Y(n4703) );
  MXI2XL U745 ( .A(n5942), .B(n3701), .S0(n366), .Y(n4702) );
  MXI2XL U746 ( .A(n5941), .B(n3700), .S0(n366), .Y(n4701) );
  MXI2XL U747 ( .A(n5940), .B(n3699), .S0(n366), .Y(n4700) );
  MXI2XL U748 ( .A(n5939), .B(n3698), .S0(n366), .Y(n4699) );
  MXI2XL U749 ( .A(n5938), .B(n3697), .S0(n366), .Y(n4698) );
  MXI2XL U750 ( .A(n5937), .B(n3696), .S0(n366), .Y(n4697) );
  MXI2XL U751 ( .A(n5936), .B(n3695), .S0(n366), .Y(n4696) );
  MXI2XL U752 ( .A(n5935), .B(n3694), .S0(n366), .Y(n4695) );
  MXI2XL U753 ( .A(n5934), .B(n3693), .S0(n366), .Y(n4694) );
  MXI2XL U754 ( .A(n5933), .B(n3692), .S0(n366), .Y(n4693) );
  MXI2XL U755 ( .A(n5932), .B(n3691), .S0(n366), .Y(n4692) );
  MXI2XL U756 ( .A(n5931), .B(n3690), .S0(n367), .Y(n4691) );
  MXI2XL U757 ( .A(n5930), .B(n3689), .S0(n367), .Y(n4690) );
  MXI2XL U758 ( .A(n5929), .B(n3688), .S0(n367), .Y(n4689) );
  MXI2XL U759 ( .A(n5928), .B(n3687), .S0(n367), .Y(n4688) );
  MXI2XL U760 ( .A(n5927), .B(n3686), .S0(n367), .Y(n4687) );
  MXI2XL U761 ( .A(n5926), .B(n3685), .S0(n367), .Y(n4686) );
  MXI2XL U762 ( .A(n5925), .B(n3684), .S0(n367), .Y(n4685) );
  MXI2XL U763 ( .A(n5924), .B(n3683), .S0(n367), .Y(n4684) );
  MXI2XL U764 ( .A(n5923), .B(n3682), .S0(n367), .Y(n4683) );
  MXI2XL U765 ( .A(n5922), .B(n3681), .S0(n367), .Y(n4682) );
  MXI2XL U766 ( .A(n5921), .B(n3680), .S0(n367), .Y(n4681) );
  MXI2XL U767 ( .A(n5920), .B(n3679), .S0(n367), .Y(n4680) );
  MXI2XL U768 ( .A(n5919), .B(n3678), .S0(n367), .Y(n4679) );
  MXI2XL U769 ( .A(n5918), .B(n3677), .S0(n368), .Y(n4678) );
  MXI2XL U770 ( .A(n5917), .B(n3676), .S0(n368), .Y(n4677) );
  MXI2XL U771 ( .A(n5916), .B(n3675), .S0(n368), .Y(n4676) );
  MXI2XL U772 ( .A(n5915), .B(n3674), .S0(n368), .Y(n4675) );
  MXI2XL U773 ( .A(n5914), .B(n3673), .S0(n368), .Y(n4674) );
  MXI2XL U774 ( .A(n5913), .B(n3672), .S0(n368), .Y(n4673) );
  MXI2XL U775 ( .A(n5912), .B(n3671), .S0(n368), .Y(n4672) );
  MXI2XL U776 ( .A(n5911), .B(n3670), .S0(n368), .Y(n4671) );
  MXI2XL U777 ( .A(n5910), .B(n3669), .S0(n368), .Y(n4670) );
  MXI2XL U778 ( .A(n5909), .B(n3668), .S0(n368), .Y(n4669) );
  MXI2XL U779 ( .A(n5908), .B(n3667), .S0(n368), .Y(n4668) );
  MXI2XL U780 ( .A(n5907), .B(n3666), .S0(n368), .Y(n4667) );
  MXI2XL U781 ( .A(n5874), .B(n3633), .S0(n3734), .Y(n4634) );
  MXI2XL U782 ( .A(n5873), .B(n3632), .S0(n366), .Y(n4633) );
  MXI2XL U783 ( .A(n5872), .B(n3631), .S0(n370), .Y(n4632) );
  MXI2XL U784 ( .A(n5871), .B(n3630), .S0(n367), .Y(n4631) );
  MXI2XL U785 ( .A(n5870), .B(n3629), .S0(n371), .Y(n4630) );
  MXI2XL U786 ( .A(n5869), .B(n3628), .S0(n364), .Y(n4629) );
  MXI2XL U787 ( .A(n5868), .B(n3627), .S0(n365), .Y(n4628) );
  MXI2XL U788 ( .A(n5867), .B(n3626), .S0(n368), .Y(n4627) );
  MXI2XL U789 ( .A(n5866), .B(n3625), .S0(n371), .Y(n4626) );
  MXI2XL U790 ( .A(n5865), .B(n3624), .S0(n371), .Y(n4625) );
  MXI2XL U791 ( .A(n5864), .B(n3623), .S0(n371), .Y(n4624) );
  MXI2XL U792 ( .A(n5863), .B(n3622), .S0(n371), .Y(n4623) );
  MXI2XL U793 ( .A(n5862), .B(n3621), .S0(n371), .Y(n4622) );
  MXI2XL U794 ( .A(n5861), .B(n3620), .S0(n371), .Y(n4621) );
  MXI2XL U795 ( .A(n5860), .B(n3619), .S0(n371), .Y(n4620) );
  MXI2XL U796 ( .A(n5859), .B(n3618), .S0(n371), .Y(n4619) );
  MXI2XL U797 ( .A(n5858), .B(n3617), .S0(n371), .Y(n4618) );
  MXI2XL U798 ( .A(n5857), .B(n3616), .S0(n371), .Y(n4617) );
  MXI2XL U799 ( .A(n5856), .B(n3615), .S0(n371), .Y(n4616) );
  MXI2XL U800 ( .A(n5855), .B(n3614), .S0(n371), .Y(n4615) );
  MXI2XL U801 ( .A(n5854), .B(n3613), .S0(n371), .Y(n4614) );
  MXI2XL U802 ( .A(n5853), .B(n3612), .S0(n365), .Y(n4613) );
  MXI2XL U803 ( .A(n5852), .B(n3611), .S0(n368), .Y(n4612) );
  MXI2XL U804 ( .A(n5851), .B(n3610), .S0(n372), .Y(n4611) );
  MXI2XL U805 ( .A(n5850), .B(n3609), .S0(n3734), .Y(n4610) );
  MXI2XL U806 ( .A(n5849), .B(n3608), .S0(n369), .Y(n4609) );
  MXI2XL U807 ( .A(n5848), .B(n3607), .S0(n366), .Y(n4608) );
  MXI2XL U808 ( .A(n5847), .B(n3606), .S0(n370), .Y(n4607) );
  MXI2XL U809 ( .A(n5846), .B(n3605), .S0(n367), .Y(n4606) );
  MXI2XL U810 ( .A(n5845), .B(n3604), .S0(n371), .Y(n4605) );
  MXI2XL U811 ( .A(n5844), .B(n3603), .S0(n364), .Y(n4604) );
  MXI2XL U812 ( .A(n5843), .B(n3602), .S0(n365), .Y(n4603) );
  MXI2XL U813 ( .A(n5815), .B(n3729), .S0(n355), .Y(n4575) );
  MXI2XL U814 ( .A(n5814), .B(n3728), .S0(n355), .Y(n4574) );
  MXI2XL U815 ( .A(n5813), .B(n3727), .S0(n355), .Y(n4573) );
  MXI2XL U816 ( .A(n5812), .B(n3726), .S0(n355), .Y(n4572) );
  MXI2XL U817 ( .A(n5811), .B(n3725), .S0(n355), .Y(n4571) );
  MXI2XL U818 ( .A(n5810), .B(n3724), .S0(n355), .Y(n4570) );
  MXI2XL U819 ( .A(n5809), .B(n3723), .S0(n355), .Y(n4569) );
  MXI2XL U820 ( .A(n5808), .B(n3722), .S0(n355), .Y(n4568) );
  MXI2XL U821 ( .A(n5807), .B(n3721), .S0(n355), .Y(n4567) );
  MXI2XL U822 ( .A(n5806), .B(n3720), .S0(n355), .Y(n4566) );
  MXI2XL U823 ( .A(n5805), .B(n3719), .S0(n355), .Y(n4565) );
  MXI2XL U824 ( .A(n5804), .B(n3718), .S0(n355), .Y(n4564) );
  MXI2XL U825 ( .A(n5803), .B(n3717), .S0(n355), .Y(n4563) );
  MXI2XL U826 ( .A(n5802), .B(n3716), .S0(n356), .Y(n4562) );
  MXI2XL U827 ( .A(n5801), .B(n3715), .S0(n356), .Y(n4561) );
  MXI2XL U828 ( .A(n5800), .B(n3714), .S0(n356), .Y(n4560) );
  MXI2XL U829 ( .A(n5799), .B(n3713), .S0(n356), .Y(n4559) );
  MXI2XL U830 ( .A(n5798), .B(n3712), .S0(n356), .Y(n4558) );
  MXI2XL U831 ( .A(n5797), .B(n3711), .S0(n356), .Y(n4557) );
  MXI2XL U832 ( .A(n5796), .B(n3710), .S0(n356), .Y(n4556) );
  MXI2XL U833 ( .A(n5795), .B(n3709), .S0(n356), .Y(n4555) );
  MXI2XL U834 ( .A(n5794), .B(n3708), .S0(n356), .Y(n4554) );
  MXI2XL U835 ( .A(n5793), .B(n3707), .S0(n356), .Y(n4553) );
  MXI2XL U836 ( .A(n5792), .B(n3706), .S0(n356), .Y(n4552) );
  MXI2XL U837 ( .A(n5791), .B(n3705), .S0(n356), .Y(n4551) );
  MXI2XL U838 ( .A(n5790), .B(n3704), .S0(n356), .Y(n4550) );
  MXI2XL U839 ( .A(n5789), .B(n3703), .S0(n357), .Y(n4549) );
  MXI2XL U840 ( .A(n5788), .B(n3702), .S0(n357), .Y(n4548) );
  MXI2XL U841 ( .A(n5787), .B(n3701), .S0(n357), .Y(n4547) );
  MXI2XL U842 ( .A(n5786), .B(n3700), .S0(n357), .Y(n4546) );
  MXI2XL U843 ( .A(n5785), .B(n3699), .S0(n357), .Y(n4545) );
  MXI2XL U844 ( .A(n5784), .B(n3698), .S0(n357), .Y(n4544) );
  MXI2XL U845 ( .A(n5783), .B(n3697), .S0(n357), .Y(n4543) );
  MXI2XL U846 ( .A(n5782), .B(n3696), .S0(n357), .Y(n4542) );
  MXI2XL U847 ( .A(n5781), .B(n3695), .S0(n357), .Y(n4541) );
  MXI2XL U848 ( .A(n5780), .B(n3694), .S0(n357), .Y(n4540) );
  MXI2XL U849 ( .A(n5779), .B(n3693), .S0(n357), .Y(n4539) );
  MXI2XL U850 ( .A(n5778), .B(n3692), .S0(n357), .Y(n4538) );
  MXI2XL U851 ( .A(n5777), .B(n3691), .S0(n357), .Y(n4537) );
  MXI2XL U852 ( .A(n5776), .B(n3690), .S0(n358), .Y(n4536) );
  MXI2XL U853 ( .A(n5775), .B(n3689), .S0(n358), .Y(n4535) );
  MXI2XL U854 ( .A(n5774), .B(n3688), .S0(n358), .Y(n4534) );
  MXI2XL U855 ( .A(n5773), .B(n3687), .S0(n358), .Y(n4533) );
  MXI2XL U856 ( .A(n5772), .B(n3686), .S0(n358), .Y(n4532) );
  MXI2XL U857 ( .A(n5771), .B(n3685), .S0(n358), .Y(n4531) );
  MXI2XL U858 ( .A(n5770), .B(n3684), .S0(n358), .Y(n4530) );
  MXI2XL U859 ( .A(n5769), .B(n3683), .S0(n358), .Y(n4529) );
  MXI2XL U860 ( .A(n5768), .B(n3682), .S0(n358), .Y(n4528) );
  MXI2XL U861 ( .A(n5767), .B(n3681), .S0(n358), .Y(n4527) );
  MXI2XL U862 ( .A(n5766), .B(n3680), .S0(n358), .Y(n4526) );
  MXI2XL U863 ( .A(n5765), .B(n3679), .S0(n358), .Y(n4525) );
  MXI2XL U864 ( .A(n5764), .B(n3678), .S0(n358), .Y(n4524) );
  MXI2XL U865 ( .A(n5763), .B(n3677), .S0(n359), .Y(n4523) );
  MXI2XL U866 ( .A(n5762), .B(n3676), .S0(n359), .Y(n4522) );
  MXI2XL U867 ( .A(n5761), .B(n3675), .S0(n359), .Y(n4521) );
  MXI2XL U868 ( .A(n5760), .B(n3674), .S0(n359), .Y(n4520) );
  MXI2XL U869 ( .A(n5759), .B(n3673), .S0(n359), .Y(n4519) );
  MXI2XL U870 ( .A(n5758), .B(n3672), .S0(n359), .Y(n4518) );
  MXI2XL U871 ( .A(n5757), .B(n3671), .S0(n359), .Y(n4517) );
  MXI2XL U872 ( .A(n5756), .B(n3670), .S0(n359), .Y(n4516) );
  MXI2XL U873 ( .A(n5755), .B(n3669), .S0(n359), .Y(n4515) );
  MXI2XL U874 ( .A(n5754), .B(n3668), .S0(n359), .Y(n4514) );
  MXI2XL U875 ( .A(n5753), .B(n3667), .S0(n359), .Y(n4513) );
  MXI2XL U876 ( .A(n5752), .B(n3666), .S0(n359), .Y(n4512) );
  MXI2XL U877 ( .A(n5719), .B(n3633), .S0(n3733), .Y(n4479) );
  MXI2XL U878 ( .A(n5718), .B(n3632), .S0(n357), .Y(n4478) );
  MXI2XL U879 ( .A(n5717), .B(n3631), .S0(n361), .Y(n4477) );
  MXI2XL U880 ( .A(n5716), .B(n3630), .S0(n358), .Y(n4476) );
  MXI2XL U881 ( .A(n5715), .B(n3629), .S0(n362), .Y(n4475) );
  MXI2XL U882 ( .A(n5714), .B(n3628), .S0(n355), .Y(n4474) );
  MXI2XL U883 ( .A(n5713), .B(n3627), .S0(n356), .Y(n4473) );
  MXI2XL U884 ( .A(n5712), .B(n3626), .S0(n359), .Y(n4472) );
  MXI2XL U885 ( .A(n5711), .B(n3625), .S0(n362), .Y(n4471) );
  MXI2XL U886 ( .A(n5710), .B(n3624), .S0(n362), .Y(n4470) );
  MXI2XL U887 ( .A(n5709), .B(n3623), .S0(n362), .Y(n4469) );
  MXI2XL U888 ( .A(n5708), .B(n3622), .S0(n362), .Y(n4468) );
  MXI2XL U889 ( .A(n5707), .B(n3621), .S0(n362), .Y(n4467) );
  MXI2XL U890 ( .A(n5706), .B(n3620), .S0(n362), .Y(n4466) );
  MXI2XL U891 ( .A(n5705), .B(n3619), .S0(n362), .Y(n4465) );
  MXI2XL U892 ( .A(n5704), .B(n3618), .S0(n362), .Y(n4464) );
  MXI2XL U893 ( .A(n5703), .B(n3617), .S0(n362), .Y(n4463) );
  MXI2XL U894 ( .A(n5702), .B(n3616), .S0(n362), .Y(n4462) );
  MXI2XL U895 ( .A(n5701), .B(n3615), .S0(n362), .Y(n4461) );
  MXI2XL U896 ( .A(n5700), .B(n3614), .S0(n362), .Y(n4460) );
  MXI2XL U897 ( .A(n5699), .B(n3613), .S0(n362), .Y(n4459) );
  MXI2XL U898 ( .A(n5698), .B(n3612), .S0(n356), .Y(n4458) );
  MXI2XL U899 ( .A(n5697), .B(n3611), .S0(n359), .Y(n4457) );
  MXI2XL U900 ( .A(n5696), .B(n3610), .S0(n363), .Y(n4456) );
  MXI2XL U901 ( .A(n5695), .B(n3609), .S0(n3733), .Y(n4455) );
  MXI2XL U902 ( .A(n5694), .B(n3608), .S0(n360), .Y(n4454) );
  MXI2XL U903 ( .A(n5693), .B(n3607), .S0(n357), .Y(n4453) );
  MXI2XL U904 ( .A(n5692), .B(n3606), .S0(n361), .Y(n4452) );
  MXI2XL U905 ( .A(n5691), .B(n3605), .S0(n358), .Y(n4451) );
  MXI2XL U906 ( .A(n5690), .B(n3604), .S0(n362), .Y(n4450) );
  MXI2XL U907 ( .A(n5689), .B(n3603), .S0(n355), .Y(n4449) );
  MXI2XL U908 ( .A(n5688), .B(n3602), .S0(n356), .Y(n4448) );
  MXI2XL U909 ( .A(n5660), .B(n3729), .S0(n345), .Y(n4420) );
  MXI2XL U910 ( .A(n5659), .B(n3728), .S0(n345), .Y(n4419) );
  MXI2XL U911 ( .A(n5658), .B(n3727), .S0(n345), .Y(n4418) );
  MXI2XL U912 ( .A(n5657), .B(n3726), .S0(n345), .Y(n4417) );
  MXI2XL U913 ( .A(n5656), .B(n3725), .S0(n345), .Y(n4416) );
  MXI2XL U914 ( .A(n5655), .B(n3724), .S0(n345), .Y(n4415) );
  MXI2XL U915 ( .A(n5654), .B(n3723), .S0(n345), .Y(n4414) );
  MXI2XL U916 ( .A(n5653), .B(n3722), .S0(n345), .Y(n4413) );
  MXI2XL U917 ( .A(n5652), .B(n3721), .S0(n345), .Y(n4412) );
  MXI2XL U918 ( .A(n5651), .B(n3720), .S0(n345), .Y(n4411) );
  MXI2XL U919 ( .A(n5650), .B(n3719), .S0(n345), .Y(n4410) );
  MXI2XL U920 ( .A(n5649), .B(n3718), .S0(n345), .Y(n4409) );
  MXI2XL U921 ( .A(n5648), .B(n3717), .S0(n345), .Y(n4408) );
  MXI2XL U922 ( .A(n5647), .B(n3716), .S0(n346), .Y(n4407) );
  MXI2XL U923 ( .A(n5646), .B(n3715), .S0(n346), .Y(n4406) );
  MXI2XL U924 ( .A(n5645), .B(n3714), .S0(n346), .Y(n4405) );
  MXI2XL U925 ( .A(n5644), .B(n3713), .S0(n346), .Y(n4404) );
  MXI2XL U926 ( .A(n5643), .B(n3712), .S0(n346), .Y(n4403) );
  MXI2XL U927 ( .A(n5642), .B(n3711), .S0(n346), .Y(n4402) );
  MXI2XL U928 ( .A(n5641), .B(n3710), .S0(n346), .Y(n4401) );
  MXI2XL U929 ( .A(n5640), .B(n3709), .S0(n346), .Y(n4400) );
  MXI2XL U930 ( .A(n5639), .B(n3708), .S0(n346), .Y(n4399) );
  MXI2XL U931 ( .A(n5638), .B(n3707), .S0(n346), .Y(n4398) );
  MXI2XL U932 ( .A(n5637), .B(n3706), .S0(n346), .Y(n4397) );
  MXI2XL U933 ( .A(n5636), .B(n3705), .S0(n346), .Y(n4396) );
  MXI2XL U934 ( .A(n5635), .B(n3704), .S0(n346), .Y(n4395) );
  MXI2XL U935 ( .A(n5634), .B(n3703), .S0(n347), .Y(n4394) );
  MXI2XL U936 ( .A(n5633), .B(n3702), .S0(n347), .Y(n4393) );
  MXI2XL U937 ( .A(n5632), .B(n3701), .S0(n347), .Y(n4392) );
  MXI2XL U938 ( .A(n5631), .B(n3700), .S0(n347), .Y(n4391) );
  MXI2XL U939 ( .A(n5630), .B(n3699), .S0(n347), .Y(n4390) );
  MXI2XL U940 ( .A(n5629), .B(n3698), .S0(n347), .Y(n4389) );
  MXI2XL U941 ( .A(n5628), .B(n3697), .S0(n347), .Y(n4388) );
  MXI2XL U942 ( .A(n5627), .B(n3696), .S0(n347), .Y(n4387) );
  MXI2XL U943 ( .A(n5626), .B(n3695), .S0(n347), .Y(n4386) );
  MXI2XL U944 ( .A(n5625), .B(n3694), .S0(n347), .Y(n4385) );
  MXI2XL U945 ( .A(n5624), .B(n3693), .S0(n347), .Y(n4384) );
  MXI2XL U946 ( .A(n5623), .B(n3692), .S0(n347), .Y(n4383) );
  MXI2XL U947 ( .A(n5622), .B(n3691), .S0(n347), .Y(n4382) );
  MXI2XL U948 ( .A(n5621), .B(n3690), .S0(n348), .Y(n4381) );
  MXI2XL U949 ( .A(n5620), .B(n3689), .S0(n348), .Y(n4380) );
  MXI2XL U950 ( .A(n5619), .B(n3688), .S0(n348), .Y(n4379) );
  MXI2XL U951 ( .A(n5618), .B(n3687), .S0(n348), .Y(n4378) );
  MXI2XL U952 ( .A(n5617), .B(n3686), .S0(n348), .Y(n4377) );
  MXI2XL U953 ( .A(n5616), .B(n3685), .S0(n348), .Y(n4376) );
  MXI2XL U954 ( .A(n5615), .B(n3684), .S0(n348), .Y(n4375) );
  MXI2XL U955 ( .A(n5614), .B(n3683), .S0(n348), .Y(n4374) );
  MXI2XL U956 ( .A(n5613), .B(n3682), .S0(n348), .Y(n4373) );
  MXI2XL U957 ( .A(n5612), .B(n3681), .S0(n348), .Y(n4372) );
  MXI2XL U958 ( .A(n5611), .B(n3680), .S0(n348), .Y(n4371) );
  MXI2XL U959 ( .A(n5610), .B(n3679), .S0(n348), .Y(n4370) );
  MXI2XL U960 ( .A(n5609), .B(n3678), .S0(n348), .Y(n4369) );
  MXI2XL U961 ( .A(n5608), .B(n3677), .S0(n349), .Y(n4368) );
  MXI2XL U962 ( .A(n5607), .B(n3676), .S0(n349), .Y(n4367) );
  MXI2XL U963 ( .A(n5606), .B(n3675), .S0(n349), .Y(n4366) );
  MXI2XL U964 ( .A(n5605), .B(n3674), .S0(n349), .Y(n4365) );
  MXI2XL U965 ( .A(n5604), .B(n3673), .S0(n349), .Y(n4364) );
  MXI2XL U966 ( .A(n5603), .B(n3672), .S0(n349), .Y(n4363) );
  MXI2XL U967 ( .A(n5602), .B(n3671), .S0(n349), .Y(n4362) );
  MXI2XL U968 ( .A(n5601), .B(n3670), .S0(n349), .Y(n4361) );
  MXI2XL U969 ( .A(n5600), .B(n3669), .S0(n349), .Y(n4360) );
  MXI2XL U970 ( .A(n5599), .B(n3668), .S0(n349), .Y(n4359) );
  MXI2XL U971 ( .A(n5598), .B(n3667), .S0(n349), .Y(n4358) );
  MXI2XL U972 ( .A(n5597), .B(n3666), .S0(n349), .Y(n4357) );
  MXI2XL U973 ( .A(n5564), .B(n3633), .S0(n3732), .Y(n4324) );
  MXI2XL U974 ( .A(n5563), .B(n3632), .S0(n347), .Y(n4323) );
  MXI2XL U975 ( .A(n5562), .B(n3631), .S0(n351), .Y(n4322) );
  MXI2XL U976 ( .A(n5561), .B(n3630), .S0(n348), .Y(n4321) );
  MXI2XL U977 ( .A(n5560), .B(n3629), .S0(n352), .Y(n4320) );
  MXI2XL U978 ( .A(n5559), .B(n3628), .S0(n345), .Y(n4319) );
  MXI2XL U979 ( .A(n5558), .B(n3627), .S0(n346), .Y(n4318) );
  MXI2XL U980 ( .A(n5557), .B(n3626), .S0(n349), .Y(n4317) );
  MXI2XL U981 ( .A(n5556), .B(n3625), .S0(n352), .Y(n4316) );
  MXI2XL U982 ( .A(n5555), .B(n3624), .S0(n352), .Y(n4315) );
  MXI2XL U983 ( .A(n5554), .B(n3623), .S0(n352), .Y(n4314) );
  MXI2XL U984 ( .A(n5553), .B(n3622), .S0(n352), .Y(n4313) );
  MXI2XL U985 ( .A(n5552), .B(n3621), .S0(n352), .Y(n4312) );
  MXI2XL U986 ( .A(n5551), .B(n3620), .S0(n352), .Y(n4311) );
  MXI2XL U987 ( .A(n5550), .B(n3619), .S0(n352), .Y(n4310) );
  MXI2XL U988 ( .A(n5549), .B(n3618), .S0(n352), .Y(n4309) );
  MXI2XL U989 ( .A(n5548), .B(n3617), .S0(n352), .Y(n4308) );
  MXI2XL U990 ( .A(n5547), .B(n3616), .S0(n352), .Y(n4307) );
  MXI2XL U991 ( .A(n5546), .B(n3615), .S0(n352), .Y(n4306) );
  MXI2XL U992 ( .A(n5545), .B(n3614), .S0(n352), .Y(n4305) );
  MXI2XL U993 ( .A(n5544), .B(n3613), .S0(n352), .Y(n4304) );
  MXI2XL U994 ( .A(n5543), .B(n3612), .S0(n346), .Y(n4303) );
  MXI2XL U995 ( .A(n5542), .B(n3611), .S0(n349), .Y(n4302) );
  MXI2XL U996 ( .A(n5541), .B(n3610), .S0(n354), .Y(n4301) );
  MXI2XL U997 ( .A(n5540), .B(n3609), .S0(n353), .Y(n4300) );
  MXI2XL U998 ( .A(n5539), .B(n3608), .S0(n350), .Y(n4299) );
  MXI2XL U999 ( .A(n5538), .B(n3607), .S0(n347), .Y(n4298) );
  MXI2XL U1000 ( .A(n5537), .B(n3606), .S0(n351), .Y(n4297) );
  MXI2XL U1001 ( .A(n5536), .B(n3605), .S0(n348), .Y(n4296) );
  MXI2XL U1002 ( .A(n5535), .B(n3604), .S0(n352), .Y(n4295) );
  MXI2XL U1003 ( .A(n5534), .B(n3603), .S0(n345), .Y(n4294) );
  MXI2XL U1004 ( .A(n5533), .B(n3602), .S0(n346), .Y(n4293) );
  MXI2XL U1005 ( .A(n5505), .B(n3729), .S0(n336), .Y(n4265) );
  MXI2XL U1006 ( .A(n5504), .B(n3728), .S0(n336), .Y(n4264) );
  MXI2XL U1007 ( .A(n5503), .B(n3727), .S0(n336), .Y(n4263) );
  MXI2XL U1008 ( .A(n5502), .B(n3726), .S0(n336), .Y(n4262) );
  MXI2XL U1009 ( .A(n5501), .B(n3725), .S0(n336), .Y(n4261) );
  MXI2XL U1010 ( .A(n5500), .B(n3724), .S0(n336), .Y(n4260) );
  MXI2XL U1011 ( .A(n5499), .B(n3723), .S0(n336), .Y(n4259) );
  MXI2XL U1012 ( .A(n5498), .B(n3722), .S0(n336), .Y(n4258) );
  MXI2XL U1013 ( .A(n5497), .B(n3721), .S0(n336), .Y(n4257) );
  MXI2XL U1014 ( .A(n5496), .B(n3720), .S0(n336), .Y(n4256) );
  MXI2XL U1015 ( .A(n5495), .B(n3719), .S0(n336), .Y(n4255) );
  MXI2XL U1016 ( .A(n5494), .B(n3718), .S0(n336), .Y(n4254) );
  MXI2XL U1017 ( .A(n5493), .B(n3717), .S0(n336), .Y(n4253) );
  MXI2XL U1018 ( .A(n5492), .B(n3716), .S0(n337), .Y(n4252) );
  MXI2XL U1019 ( .A(n5491), .B(n3715), .S0(n337), .Y(n4251) );
  MXI2XL U1020 ( .A(n5490), .B(n3714), .S0(n337), .Y(n4250) );
  MXI2XL U1021 ( .A(n5489), .B(n3713), .S0(n337), .Y(n4249) );
  MXI2XL U1022 ( .A(n5488), .B(n3712), .S0(n337), .Y(n4248) );
  MXI2XL U1023 ( .A(n5487), .B(n3711), .S0(n337), .Y(n4247) );
  MXI2XL U1024 ( .A(n5486), .B(n3710), .S0(n337), .Y(n4246) );
  MXI2XL U1025 ( .A(n5485), .B(n3709), .S0(n337), .Y(n4245) );
  MXI2XL U1026 ( .A(n5484), .B(n3708), .S0(n337), .Y(n4244) );
  MXI2XL U1027 ( .A(n5483), .B(n3707), .S0(n337), .Y(n4243) );
  MXI2XL U1028 ( .A(n5482), .B(n3706), .S0(n337), .Y(n4242) );
  MXI2XL U1029 ( .A(n5481), .B(n3705), .S0(n337), .Y(n4241) );
  MXI2XL U1030 ( .A(n5480), .B(n3704), .S0(n337), .Y(n4240) );
  MXI2XL U1031 ( .A(n5479), .B(n3703), .S0(n338), .Y(n4239) );
  MXI2XL U1032 ( .A(n5478), .B(n3702), .S0(n338), .Y(n4238) );
  MXI2XL U1033 ( .A(n5477), .B(n3701), .S0(n338), .Y(n4237) );
  MXI2XL U1034 ( .A(n5476), .B(n3700), .S0(n338), .Y(n4236) );
  MXI2XL U1035 ( .A(n5475), .B(n3699), .S0(n338), .Y(n4235) );
  MXI2XL U1036 ( .A(n5474), .B(n3698), .S0(n338), .Y(n4234) );
  MXI2XL U1037 ( .A(n5473), .B(n3697), .S0(n338), .Y(n4233) );
  MXI2XL U1038 ( .A(n5472), .B(n3696), .S0(n338), .Y(n4232) );
  MXI2XL U1039 ( .A(n5471), .B(n3695), .S0(n338), .Y(n4231) );
  MXI2XL U1040 ( .A(n5470), .B(n3694), .S0(n338), .Y(n4230) );
  MXI2XL U1041 ( .A(n5469), .B(n3693), .S0(n338), .Y(n4229) );
  MXI2XL U1042 ( .A(n5468), .B(n3692), .S0(n338), .Y(n4228) );
  MXI2XL U1043 ( .A(n5467), .B(n3691), .S0(n338), .Y(n4227) );
  MXI2XL U1044 ( .A(n5466), .B(n3690), .S0(n339), .Y(n4226) );
  MXI2XL U1045 ( .A(n5465), .B(n3689), .S0(n339), .Y(n4225) );
  MXI2XL U1046 ( .A(n5464), .B(n3688), .S0(n339), .Y(n4224) );
  MXI2XL U1047 ( .A(n5463), .B(n3687), .S0(n339), .Y(n4223) );
  MXI2XL U1048 ( .A(n5462), .B(n3686), .S0(n339), .Y(n4222) );
  MXI2XL U1049 ( .A(n5461), .B(n3685), .S0(n339), .Y(n4221) );
  MXI2XL U1050 ( .A(n5460), .B(n3684), .S0(n339), .Y(n4220) );
  MXI2XL U1051 ( .A(n5459), .B(n3683), .S0(n339), .Y(n4219) );
  MXI2XL U1052 ( .A(n5458), .B(n3682), .S0(n339), .Y(n4218) );
  MXI2XL U1053 ( .A(n5457), .B(n3681), .S0(n339), .Y(n4217) );
  MXI2XL U1054 ( .A(n5456), .B(n3680), .S0(n339), .Y(n4216) );
  MXI2XL U1055 ( .A(n5455), .B(n3679), .S0(n339), .Y(n4215) );
  MXI2XL U1056 ( .A(n5454), .B(n3678), .S0(n339), .Y(n4214) );
  MXI2XL U1057 ( .A(n5453), .B(n3677), .S0(n340), .Y(n4213) );
  MXI2XL U1058 ( .A(n5452), .B(n3676), .S0(n340), .Y(n4212) );
  MXI2XL U1059 ( .A(n5451), .B(n3675), .S0(n340), .Y(n4211) );
  MXI2XL U1060 ( .A(n5450), .B(n3674), .S0(n340), .Y(n4210) );
  MXI2XL U1061 ( .A(n5449), .B(n3673), .S0(n340), .Y(n4209) );
  MXI2XL U1062 ( .A(n5448), .B(n3672), .S0(n340), .Y(n4208) );
  MXI2XL U1063 ( .A(n5447), .B(n3671), .S0(n340), .Y(n4207) );
  MXI2XL U1064 ( .A(n5446), .B(n3670), .S0(n340), .Y(n4206) );
  MXI2XL U1065 ( .A(n5445), .B(n3669), .S0(n340), .Y(n4205) );
  MXI2XL U1066 ( .A(n5444), .B(n3668), .S0(n340), .Y(n4204) );
  MXI2XL U1067 ( .A(n5443), .B(n3667), .S0(n340), .Y(n4203) );
  MXI2XL U1068 ( .A(n5442), .B(n3666), .S0(n340), .Y(n4202) );
  MXI2XL U1069 ( .A(n5409), .B(n3633), .S0(n3731), .Y(n4169) );
  MXI2XL U1070 ( .A(n5408), .B(n3632), .S0(n338), .Y(n4168) );
  MXI2XL U1071 ( .A(n5407), .B(n3631), .S0(n342), .Y(n4167) );
  MXI2XL U1072 ( .A(n5406), .B(n3630), .S0(n339), .Y(n4166) );
  MXI2XL U1073 ( .A(n5405), .B(n3629), .S0(n343), .Y(n4165) );
  MXI2XL U1074 ( .A(n5404), .B(n3628), .S0(n336), .Y(n4164) );
  MXI2XL U1075 ( .A(n5403), .B(n3627), .S0(n337), .Y(n4163) );
  MXI2XL U1076 ( .A(n5402), .B(n3626), .S0(n340), .Y(n4162) );
  MXI2XL U1077 ( .A(n5401), .B(n3625), .S0(n343), .Y(n4161) );
  MXI2XL U1078 ( .A(n5400), .B(n3624), .S0(n343), .Y(n4160) );
  MXI2XL U1079 ( .A(n5399), .B(n3623), .S0(n343), .Y(n4159) );
  MXI2XL U1080 ( .A(n5398), .B(n3622), .S0(n343), .Y(n4158) );
  MXI2XL U1081 ( .A(n5397), .B(n3621), .S0(n343), .Y(n4157) );
  MXI2XL U1082 ( .A(n5396), .B(n3620), .S0(n343), .Y(n4156) );
  MXI2XL U1083 ( .A(n5395), .B(n3619), .S0(n343), .Y(n4155) );
  MXI2XL U1084 ( .A(n5394), .B(n3618), .S0(n343), .Y(n4154) );
  MXI2XL U1085 ( .A(n5393), .B(n3617), .S0(n343), .Y(n4153) );
  MXI2XL U1086 ( .A(n5392), .B(n3616), .S0(n343), .Y(n4152) );
  MXI2XL U1087 ( .A(n5391), .B(n3615), .S0(n343), .Y(n4151) );
  MXI2XL U1088 ( .A(n5390), .B(n3614), .S0(n343), .Y(n4150) );
  MXI2XL U1089 ( .A(n5389), .B(n3613), .S0(n343), .Y(n4149) );
  MXI2XL U1090 ( .A(n5388), .B(n3612), .S0(n337), .Y(n4148) );
  MXI2XL U1091 ( .A(n5387), .B(n3611), .S0(n340), .Y(n4147) );
  MXI2XL U1092 ( .A(n5386), .B(n3610), .S0(n344), .Y(n4146) );
  MXI2XL U1093 ( .A(n5385), .B(n3609), .S0(n3731), .Y(n4145) );
  MXI2XL U1094 ( .A(n5384), .B(n3608), .S0(n341), .Y(n4144) );
  MXI2XL U1095 ( .A(n5383), .B(n3607), .S0(n338), .Y(n4143) );
  MXI2XL U1096 ( .A(n5382), .B(n3606), .S0(n342), .Y(n4142) );
  MXI2XL U1097 ( .A(n5381), .B(n3605), .S0(n339), .Y(n4141) );
  MXI2XL U1098 ( .A(n5380), .B(n3604), .S0(n343), .Y(n4140) );
  MXI2XL U1099 ( .A(n5379), .B(n3603), .S0(n336), .Y(n4139) );
  MXI2XL U1100 ( .A(n5378), .B(n3602), .S0(n337), .Y(n4138) );
  MXI2XL U1101 ( .A(n5350), .B(n3729), .S0(n327), .Y(n4110) );
  MXI2XL U1102 ( .A(n5349), .B(n3728), .S0(n327), .Y(n4109) );
  MXI2XL U1103 ( .A(n5348), .B(n3727), .S0(n327), .Y(n4108) );
  MXI2XL U1104 ( .A(n5347), .B(n3726), .S0(n327), .Y(n4107) );
  MXI2XL U1105 ( .A(n5346), .B(n3725), .S0(n327), .Y(n4106) );
  MXI2XL U1106 ( .A(n5345), .B(n3724), .S0(n327), .Y(n4105) );
  MXI2XL U1107 ( .A(n5344), .B(n3723), .S0(n327), .Y(n4104) );
  MXI2XL U1108 ( .A(n5343), .B(n3722), .S0(n327), .Y(n4103) );
  MXI2XL U1109 ( .A(n5342), .B(n3721), .S0(n327), .Y(n4102) );
  MXI2XL U1110 ( .A(n5341), .B(n3720), .S0(n327), .Y(n4101) );
  MXI2XL U1111 ( .A(n5340), .B(n3719), .S0(n327), .Y(n4100) );
  MXI2XL U1112 ( .A(n5339), .B(n3718), .S0(n327), .Y(n4099) );
  MXI2XL U1113 ( .A(n5338), .B(n3717), .S0(n327), .Y(n4098) );
  MXI2XL U1114 ( .A(n5337), .B(n3716), .S0(n328), .Y(n4097) );
  MXI2XL U1115 ( .A(n5336), .B(n3715), .S0(n328), .Y(n4096) );
  MXI2XL U1116 ( .A(n5335), .B(n3714), .S0(n328), .Y(n4095) );
  MXI2XL U1117 ( .A(n5334), .B(n3713), .S0(n328), .Y(n4094) );
  MXI2XL U1118 ( .A(n5333), .B(n3712), .S0(n328), .Y(n4093) );
  MXI2XL U1119 ( .A(n5332), .B(n3711), .S0(n328), .Y(n4092) );
  MXI2XL U1120 ( .A(n5331), .B(n3710), .S0(n328), .Y(n4091) );
  MXI2XL U1121 ( .A(n5330), .B(n3709), .S0(n328), .Y(n4090) );
  MXI2XL U1122 ( .A(n5329), .B(n3708), .S0(n328), .Y(n4089) );
  MXI2XL U1123 ( .A(n5328), .B(n3707), .S0(n328), .Y(n4088) );
  MXI2XL U1124 ( .A(n5327), .B(n3706), .S0(n328), .Y(n4087) );
  MXI2XL U1125 ( .A(n5326), .B(n3705), .S0(n328), .Y(n4086) );
  MXI2XL U1126 ( .A(n5325), .B(n3704), .S0(n328), .Y(n4085) );
  MXI2XL U1127 ( .A(n5324), .B(n3703), .S0(n329), .Y(n4084) );
  MXI2XL U1128 ( .A(n5323), .B(n3702), .S0(n329), .Y(n4083) );
  MXI2XL U1129 ( .A(n5322), .B(n3701), .S0(n329), .Y(n4082) );
  MXI2XL U1130 ( .A(n5321), .B(n3700), .S0(n329), .Y(n4081) );
  MXI2XL U1131 ( .A(n5320), .B(n3699), .S0(n329), .Y(n4080) );
  MXI2XL U1132 ( .A(n5319), .B(n3698), .S0(n329), .Y(n4079) );
  MXI2XL U1133 ( .A(n5318), .B(n3697), .S0(n329), .Y(n4078) );
  MXI2XL U1134 ( .A(n5317), .B(n3696), .S0(n329), .Y(n4077) );
  MXI2XL U1135 ( .A(n5316), .B(n3695), .S0(n329), .Y(n4076) );
  MXI2XL U1136 ( .A(n5315), .B(n3694), .S0(n329), .Y(n4075) );
  MXI2XL U1137 ( .A(n5314), .B(n3693), .S0(n329), .Y(n4074) );
  MXI2XL U1138 ( .A(n5313), .B(n3692), .S0(n329), .Y(n4073) );
  MXI2XL U1139 ( .A(n5312), .B(n3691), .S0(n329), .Y(n4072) );
  MXI2XL U1140 ( .A(n5311), .B(n3690), .S0(n330), .Y(n4071) );
  MXI2XL U1141 ( .A(n5310), .B(n3689), .S0(n330), .Y(n4070) );
  MXI2XL U1142 ( .A(n5309), .B(n3688), .S0(n330), .Y(n4069) );
  MXI2XL U1143 ( .A(n5308), .B(n3687), .S0(n330), .Y(n4068) );
  MXI2XL U1144 ( .A(n5307), .B(n3686), .S0(n330), .Y(n4067) );
  MXI2XL U1145 ( .A(n5306), .B(n3685), .S0(n330), .Y(n4066) );
  MXI2XL U1146 ( .A(n5305), .B(n3684), .S0(n330), .Y(n4065) );
  MXI2XL U1147 ( .A(n5304), .B(n3683), .S0(n330), .Y(n4064) );
  MXI2XL U1148 ( .A(n5303), .B(n3682), .S0(n330), .Y(n4063) );
  MXI2XL U1149 ( .A(n5302), .B(n3681), .S0(n330), .Y(n4062) );
  MXI2XL U1150 ( .A(n5301), .B(n3680), .S0(n330), .Y(n4061) );
  MXI2XL U1151 ( .A(n5300), .B(n3679), .S0(n330), .Y(n4060) );
  MXI2XL U1152 ( .A(n5299), .B(n3678), .S0(n330), .Y(n4059) );
  MXI2XL U1153 ( .A(n5298), .B(n3677), .S0(n331), .Y(n4058) );
  MXI2XL U1154 ( .A(n5297), .B(n3676), .S0(n331), .Y(n4057) );
  MXI2XL U1155 ( .A(n5296), .B(n3675), .S0(n331), .Y(n4056) );
  MXI2XL U1156 ( .A(n5295), .B(n3674), .S0(n331), .Y(n4055) );
  MXI2XL U1157 ( .A(n5294), .B(n3673), .S0(n331), .Y(n4054) );
  MXI2XL U1158 ( .A(n5293), .B(n3672), .S0(n331), .Y(n4053) );
  MXI2XL U1159 ( .A(n5292), .B(n3671), .S0(n331), .Y(n4052) );
  MXI2XL U1160 ( .A(n5291), .B(n3670), .S0(n331), .Y(n4051) );
  MXI2XL U1161 ( .A(n5290), .B(n3669), .S0(n331), .Y(n4050) );
  MXI2XL U1162 ( .A(n5289), .B(n3668), .S0(n331), .Y(n4049) );
  MXI2XL U1163 ( .A(n5288), .B(n3667), .S0(n331), .Y(n4048) );
  MXI2XL U1164 ( .A(n5287), .B(n3666), .S0(n331), .Y(n4047) );
  MXI2XL U1165 ( .A(n5254), .B(n3633), .S0(n3730), .Y(n4014) );
  MXI2XL U1166 ( .A(n5253), .B(n3632), .S0(n329), .Y(n4013) );
  MXI2XL U1167 ( .A(n5252), .B(n3631), .S0(n333), .Y(n4012) );
  MXI2XL U1168 ( .A(n5251), .B(n3630), .S0(n330), .Y(n4011) );
  MXI2XL U1169 ( .A(n5250), .B(n3629), .S0(n334), .Y(n4010) );
  MXI2XL U1170 ( .A(n5249), .B(n3628), .S0(n327), .Y(n4009) );
  MXI2XL U1171 ( .A(n5248), .B(n3627), .S0(n328), .Y(n4008) );
  MXI2XL U1172 ( .A(n5247), .B(n3626), .S0(n331), .Y(n4007) );
  MXI2XL U1173 ( .A(n5246), .B(n3625), .S0(n334), .Y(n4006) );
  MXI2XL U1174 ( .A(n5245), .B(n3624), .S0(n334), .Y(n4005) );
  MXI2XL U1175 ( .A(n5244), .B(n3623), .S0(n334), .Y(n4004) );
  MXI2XL U1176 ( .A(n5243), .B(n3622), .S0(n334), .Y(n4003) );
  MXI2XL U1177 ( .A(n5242), .B(n3621), .S0(n334), .Y(n4002) );
  MXI2XL U1178 ( .A(n5241), .B(n3620), .S0(n334), .Y(n4001) );
  MXI2XL U1179 ( .A(n5240), .B(n3619), .S0(n334), .Y(n4000) );
  MXI2XL U1180 ( .A(n5239), .B(n3618), .S0(n334), .Y(n3999) );
  MXI2XL U1181 ( .A(n5238), .B(n3617), .S0(n334), .Y(n3998) );
  MXI2XL U1182 ( .A(n5237), .B(n3616), .S0(n334), .Y(n3997) );
  MXI2XL U1183 ( .A(n5236), .B(n3615), .S0(n334), .Y(n3996) );
  MXI2XL U1184 ( .A(n5235), .B(n3614), .S0(n334), .Y(n3995) );
  MXI2XL U1185 ( .A(n5234), .B(n3613), .S0(n334), .Y(n3994) );
  MXI2XL U1186 ( .A(n5233), .B(n3612), .S0(n328), .Y(n3993) );
  MXI2XL U1187 ( .A(n5232), .B(n3611), .S0(n331), .Y(n3992) );
  MXI2XL U1188 ( .A(n5231), .B(n3610), .S0(n335), .Y(n3991) );
  MXI2XL U1189 ( .A(n5230), .B(n3609), .S0(n3730), .Y(n3990) );
  MXI2XL U1190 ( .A(n5229), .B(n3608), .S0(n332), .Y(n3989) );
  MXI2XL U1191 ( .A(n5228), .B(n3607), .S0(n329), .Y(n3988) );
  MXI2XL U1192 ( .A(n5227), .B(n3606), .S0(n333), .Y(n3987) );
  MXI2XL U1193 ( .A(n5226), .B(n3605), .S0(n330), .Y(n3986) );
  MXI2XL U1194 ( .A(n5225), .B(n3604), .S0(n334), .Y(n3985) );
  MXI2XL U1195 ( .A(n5224), .B(n3603), .S0(n327), .Y(n3984) );
  MXI2XL U1196 ( .A(n5223), .B(n3602), .S0(n328), .Y(n3983) );
  MXI2XL U1197 ( .A(n5195), .B(n3729), .S0(n318), .Y(n3955) );
  MXI2XL U1198 ( .A(n5194), .B(n3728), .S0(n318), .Y(n3954) );
  MXI2XL U1199 ( .A(n5193), .B(n3727), .S0(n318), .Y(n3953) );
  MXI2XL U1200 ( .A(n5192), .B(n3726), .S0(n318), .Y(n3952) );
  MXI2XL U1201 ( .A(n5191), .B(n3725), .S0(n318), .Y(n3951) );
  MXI2XL U1202 ( .A(n5190), .B(n3724), .S0(n318), .Y(n3950) );
  MXI2XL U1203 ( .A(n5189), .B(n3723), .S0(n318), .Y(n3949) );
  MXI2XL U1204 ( .A(n5188), .B(n3722), .S0(n318), .Y(n3948) );
  MXI2XL U1205 ( .A(n5187), .B(n3721), .S0(n318), .Y(n3947) );
  MXI2XL U1206 ( .A(n5186), .B(n3720), .S0(n318), .Y(n3946) );
  MXI2XL U1207 ( .A(n5185), .B(n3719), .S0(n318), .Y(n3945) );
  MXI2XL U1208 ( .A(n5184), .B(n3718), .S0(n318), .Y(n3944) );
  MXI2XL U1209 ( .A(n5183), .B(n3717), .S0(n318), .Y(n3943) );
  MXI2XL U1210 ( .A(n5182), .B(n3716), .S0(n319), .Y(n3942) );
  MXI2XL U1211 ( .A(n5181), .B(n3715), .S0(n319), .Y(n3941) );
  MXI2XL U1212 ( .A(n5180), .B(n3714), .S0(n319), .Y(n3940) );
  MXI2XL U1213 ( .A(n5179), .B(n3713), .S0(n319), .Y(n3939) );
  MXI2XL U1214 ( .A(n5178), .B(n3712), .S0(n319), .Y(n3938) );
  MXI2XL U1215 ( .A(n5177), .B(n3711), .S0(n319), .Y(n3937) );
  MXI2XL U1216 ( .A(n5176), .B(n3710), .S0(n319), .Y(n3936) );
  MXI2XL U1217 ( .A(n5175), .B(n3709), .S0(n319), .Y(n3935) );
  MXI2XL U1218 ( .A(n5174), .B(n3708), .S0(n319), .Y(n3934) );
  MXI2XL U1219 ( .A(n5173), .B(n3707), .S0(n319), .Y(n3933) );
  MXI2XL U1220 ( .A(n5172), .B(n3706), .S0(n319), .Y(n3932) );
  MXI2XL U1221 ( .A(n5171), .B(n3705), .S0(n319), .Y(n3931) );
  MXI2XL U1222 ( .A(n5170), .B(n3704), .S0(n319), .Y(n3930) );
  MXI2XL U1223 ( .A(n5169), .B(n3703), .S0(n320), .Y(n3929) );
  MXI2XL U1224 ( .A(n5168), .B(n3702), .S0(n320), .Y(n3928) );
  MXI2XL U1225 ( .A(n5167), .B(n3701), .S0(n320), .Y(n3927) );
  MXI2XL U1226 ( .A(n5166), .B(n3700), .S0(n320), .Y(n3926) );
  MXI2XL U1227 ( .A(n5165), .B(n3699), .S0(n320), .Y(n3925) );
  MXI2XL U1228 ( .A(n5164), .B(n3698), .S0(n320), .Y(n3924) );
  MXI2XL U1229 ( .A(n5163), .B(n3697), .S0(n320), .Y(n3923) );
  MXI2XL U1230 ( .A(n5162), .B(n3696), .S0(n320), .Y(n3922) );
  MXI2XL U1231 ( .A(n5161), .B(n3695), .S0(n320), .Y(n3921) );
  MXI2XL U1232 ( .A(n5160), .B(n3694), .S0(n320), .Y(n3920) );
  MXI2XL U1233 ( .A(n5159), .B(n3693), .S0(n320), .Y(n3919) );
  MXI2XL U1234 ( .A(n5158), .B(n3692), .S0(n320), .Y(n3918) );
  MXI2XL U1235 ( .A(n5157), .B(n3691), .S0(n320), .Y(n3917) );
  MXI2XL U1236 ( .A(n5156), .B(n3690), .S0(n321), .Y(n3916) );
  MXI2XL U1237 ( .A(n5155), .B(n3689), .S0(n321), .Y(n3915) );
  MXI2XL U1238 ( .A(n5154), .B(n3688), .S0(n321), .Y(n3914) );
  MXI2XL U1239 ( .A(n5153), .B(n3687), .S0(n321), .Y(n3913) );
  MXI2XL U1240 ( .A(n5152), .B(n3686), .S0(n321), .Y(n3912) );
  MXI2XL U1241 ( .A(n5151), .B(n3685), .S0(n321), .Y(n3911) );
  MXI2XL U1242 ( .A(n5150), .B(n3684), .S0(n321), .Y(n3910) );
  MXI2XL U1243 ( .A(n5149), .B(n3683), .S0(n321), .Y(n3909) );
  MXI2XL U1244 ( .A(n5148), .B(n3682), .S0(n321), .Y(n3908) );
  MXI2XL U1245 ( .A(n5147), .B(n3681), .S0(n321), .Y(n3907) );
  MXI2XL U1246 ( .A(n5146), .B(n3680), .S0(n321), .Y(n3906) );
  MXI2XL U1247 ( .A(n5145), .B(n3679), .S0(n321), .Y(n3905) );
  MXI2XL U1248 ( .A(n5144), .B(n3678), .S0(n321), .Y(n3904) );
  MXI2XL U1249 ( .A(n5143), .B(n3677), .S0(n322), .Y(n3903) );
  MXI2XL U1250 ( .A(n5142), .B(n3676), .S0(n322), .Y(n3902) );
  MXI2XL U1251 ( .A(n5141), .B(n3675), .S0(n322), .Y(n3901) );
  MXI2XL U1252 ( .A(n5140), .B(n3674), .S0(n322), .Y(n3900) );
  MXI2XL U1253 ( .A(n5139), .B(n3673), .S0(n322), .Y(n3899) );
  MXI2XL U1254 ( .A(n5138), .B(n3672), .S0(n322), .Y(n3898) );
  MXI2XL U1255 ( .A(n5137), .B(n3671), .S0(n322), .Y(n3897) );
  MXI2XL U1256 ( .A(n5136), .B(n3670), .S0(n322), .Y(n3896) );
  MXI2XL U1257 ( .A(n5135), .B(n3669), .S0(n322), .Y(n3895) );
  MXI2XL U1258 ( .A(n5134), .B(n3668), .S0(n322), .Y(n3894) );
  MXI2XL U1259 ( .A(n5133), .B(n3667), .S0(n322), .Y(n3893) );
  MXI2XL U1260 ( .A(n5132), .B(n3666), .S0(n322), .Y(n3892) );
  MXI2XL U1261 ( .A(n5099), .B(n3633), .S0(n3575), .Y(n3859) );
  MXI2XL U1262 ( .A(n5098), .B(n3632), .S0(n320), .Y(n3858) );
  MXI2XL U1263 ( .A(n5097), .B(n3631), .S0(n324), .Y(n3857) );
  MXI2XL U1264 ( .A(n5096), .B(n3630), .S0(n321), .Y(n3856) );
  MXI2XL U1265 ( .A(n5095), .B(n3629), .S0(n325), .Y(n3855) );
  MXI2XL U1266 ( .A(n5094), .B(n3628), .S0(n318), .Y(n3854) );
  MXI2XL U1267 ( .A(n5093), .B(n3627), .S0(n319), .Y(n3853) );
  MXI2XL U1268 ( .A(n5092), .B(n3626), .S0(n322), .Y(n3852) );
  MXI2XL U1269 ( .A(n5091), .B(n3625), .S0(n325), .Y(n3851) );
  MXI2XL U1270 ( .A(n5090), .B(n3624), .S0(n325), .Y(n3850) );
  MXI2XL U1271 ( .A(n5089), .B(n3623), .S0(n325), .Y(n3849) );
  MXI2XL U1272 ( .A(n5088), .B(n3622), .S0(n325), .Y(n3848) );
  MXI2XL U1273 ( .A(n5087), .B(n3621), .S0(n325), .Y(n3847) );
  MXI2XL U1274 ( .A(n5086), .B(n3620), .S0(n325), .Y(n3846) );
  MXI2XL U1275 ( .A(n5085), .B(n3619), .S0(n325), .Y(n3845) );
  MXI2XL U1276 ( .A(n5084), .B(n3618), .S0(n325), .Y(n3844) );
  MXI2XL U1277 ( .A(n5083), .B(n3617), .S0(n325), .Y(n3843) );
  MXI2XL U1278 ( .A(n5082), .B(n3616), .S0(n325), .Y(n3842) );
  MXI2XL U1279 ( .A(n5081), .B(n3615), .S0(n325), .Y(n3841) );
  MXI2XL U1280 ( .A(n5080), .B(n3614), .S0(n325), .Y(n3840) );
  MXI2XL U1281 ( .A(n5079), .B(n3613), .S0(n325), .Y(n3839) );
  MXI2XL U1282 ( .A(n5078), .B(n3612), .S0(n319), .Y(n3838) );
  MXI2XL U1283 ( .A(n5077), .B(n3611), .S0(n322), .Y(n3837) );
  MXI2XL U1284 ( .A(n5076), .B(n3610), .S0(n326), .Y(n3836) );
  MXI2XL U1285 ( .A(n5075), .B(n3609), .S0(n3575), .Y(n3835) );
  MXI2XL U1286 ( .A(n5074), .B(n3608), .S0(n323), .Y(n3834) );
  MXI2XL U1287 ( .A(n5073), .B(n3607), .S0(n320), .Y(n3833) );
  MXI2XL U1288 ( .A(n5072), .B(n3606), .S0(n324), .Y(n3832) );
  MXI2XL U1289 ( .A(n5071), .B(n3605), .S0(n321), .Y(n3831) );
  MXI2XL U1290 ( .A(n5070), .B(n3604), .S0(n325), .Y(n3830) );
  MXI2XL U1291 ( .A(n5069), .B(n3603), .S0(n318), .Y(n3829) );
  MXI2XL U1292 ( .A(n5068), .B(n3602), .S0(n319), .Y(n3828) );
  MXI2XL U1293 ( .A(n6216), .B(n3665), .S0(n386), .Y(n4976) );
  MXI2XL U1294 ( .A(n6215), .B(n3664), .S0(n387), .Y(n4975) );
  MXI2XL U1295 ( .A(n6214), .B(n3663), .S0(n387), .Y(n4974) );
  MXI2XL U1296 ( .A(n6213), .B(n3662), .S0(n387), .Y(n4973) );
  MXI2XL U1297 ( .A(n6212), .B(n3661), .S0(n387), .Y(n4972) );
  MXI2XL U1298 ( .A(n6211), .B(n3660), .S0(n387), .Y(n4971) );
  MXI2XL U1299 ( .A(n6210), .B(n3659), .S0(n387), .Y(n4970) );
  MXI2XL U1300 ( .A(n6209), .B(n3658), .S0(n387), .Y(n4969) );
  MXI2XL U1301 ( .A(n6208), .B(n3657), .S0(n387), .Y(n4968) );
  MXI2XL U1302 ( .A(n6207), .B(n3656), .S0(n387), .Y(n4967) );
  MXI2XL U1303 ( .A(n6206), .B(n3655), .S0(n387), .Y(n4966) );
  MXI2XL U1304 ( .A(n6205), .B(n3654), .S0(n387), .Y(n4965) );
  MXI2XL U1305 ( .A(n6204), .B(n3653), .S0(n387), .Y(n4964) );
  MXI2XL U1306 ( .A(n6203), .B(n3652), .S0(n387), .Y(n4963) );
  MXI2XL U1307 ( .A(n6202), .B(n3651), .S0(n388), .Y(n4962) );
  MXI2XL U1308 ( .A(n6201), .B(n3650), .S0(n388), .Y(n4961) );
  MXI2XL U1309 ( .A(n6200), .B(n3649), .S0(n388), .Y(n4960) );
  MXI2XL U1310 ( .A(n6199), .B(n3648), .S0(n388), .Y(n4959) );
  MXI2XL U1311 ( .A(n6198), .B(n3647), .S0(n388), .Y(n4958) );
  MXI2XL U1312 ( .A(n6197), .B(n3646), .S0(n388), .Y(n4957) );
  MXI2XL U1313 ( .A(n6196), .B(n3645), .S0(n388), .Y(n4956) );
  MXI2XL U1314 ( .A(n6195), .B(n3644), .S0(n388), .Y(n4955) );
  MXI2XL U1315 ( .A(n6194), .B(n3643), .S0(n388), .Y(n4954) );
  MXI2XL U1316 ( .A(n6193), .B(n3642), .S0(n388), .Y(n4953) );
  MXI2XL U1317 ( .A(n6192), .B(n3641), .S0(n388), .Y(n4952) );
  MXI2XL U1318 ( .A(n6191), .B(n3640), .S0(n388), .Y(n4951) );
  MXI2XL U1319 ( .A(n6190), .B(n3639), .S0(n388), .Y(n4950) );
  MXI2XL U1320 ( .A(n6189), .B(n3638), .S0(n382), .Y(n4949) );
  MXI2XL U1321 ( .A(n6188), .B(n3637), .S0(n384), .Y(n4948) );
  MXI2XL U1322 ( .A(n6187), .B(n3636), .S0(n388), .Y(n4947) );
  MXI2XL U1323 ( .A(n6186), .B(n3635), .S0(n385), .Y(n4946) );
  MXI2XL U1324 ( .A(n6185), .B(n3634), .S0(n389), .Y(n4945) );
  MXI2XL U1325 ( .A(n6061), .B(n3665), .S0(n377), .Y(n4821) );
  MXI2XL U1326 ( .A(n6060), .B(n3664), .S0(n378), .Y(n4820) );
  MXI2XL U1327 ( .A(n6059), .B(n3663), .S0(n378), .Y(n4819) );
  MXI2XL U1328 ( .A(n6058), .B(n3662), .S0(n378), .Y(n4818) );
  MXI2XL U1329 ( .A(n6057), .B(n3661), .S0(n378), .Y(n4817) );
  MXI2XL U1330 ( .A(n6056), .B(n3660), .S0(n378), .Y(n4816) );
  MXI2XL U1331 ( .A(n6055), .B(n3659), .S0(n378), .Y(n4815) );
  MXI2XL U1332 ( .A(n6054), .B(n3658), .S0(n378), .Y(n4814) );
  MXI2XL U1333 ( .A(n6053), .B(n3657), .S0(n378), .Y(n4813) );
  MXI2XL U1334 ( .A(n6052), .B(n3656), .S0(n378), .Y(n4812) );
  MXI2XL U1335 ( .A(n6051), .B(n3655), .S0(n378), .Y(n4811) );
  MXI2XL U1336 ( .A(n6050), .B(n3654), .S0(n378), .Y(n4810) );
  MXI2XL U1337 ( .A(n6049), .B(n3653), .S0(n378), .Y(n4809) );
  MXI2XL U1338 ( .A(n6048), .B(n3652), .S0(n378), .Y(n4808) );
  MXI2XL U1339 ( .A(n6047), .B(n3651), .S0(n379), .Y(n4807) );
  MXI2XL U1340 ( .A(n6046), .B(n3650), .S0(n379), .Y(n4806) );
  MXI2XL U1341 ( .A(n6045), .B(n3649), .S0(n379), .Y(n4805) );
  MXI2XL U1342 ( .A(n6044), .B(n3648), .S0(n379), .Y(n4804) );
  MXI2XL U1343 ( .A(n6043), .B(n3647), .S0(n379), .Y(n4803) );
  MXI2XL U1344 ( .A(n6042), .B(n3646), .S0(n379), .Y(n4802) );
  MXI2XL U1345 ( .A(n6041), .B(n3645), .S0(n379), .Y(n4801) );
  MXI2XL U1346 ( .A(n6040), .B(n3644), .S0(n379), .Y(n4800) );
  MXI2XL U1347 ( .A(n6039), .B(n3643), .S0(n379), .Y(n4799) );
  MXI2XL U1348 ( .A(n6038), .B(n3642), .S0(n379), .Y(n4798) );
  MXI2XL U1349 ( .A(n6037), .B(n3641), .S0(n379), .Y(n4797) );
  MXI2XL U1350 ( .A(n6036), .B(n3640), .S0(n379), .Y(n4796) );
  MXI2XL U1351 ( .A(n6035), .B(n3639), .S0(n379), .Y(n4795) );
  MXI2XL U1352 ( .A(n6034), .B(n3638), .S0(n373), .Y(n4794) );
  MXI2XL U1353 ( .A(n6033), .B(n3637), .S0(n375), .Y(n4793) );
  MXI2XL U1354 ( .A(n6032), .B(n3636), .S0(n379), .Y(n4792) );
  MXI2XL U1355 ( .A(n6031), .B(n3635), .S0(n376), .Y(n4791) );
  MXI2XL U1356 ( .A(n6030), .B(n3634), .S0(n380), .Y(n4790) );
  MXI2XL U1357 ( .A(n5906), .B(n3665), .S0(n368), .Y(n4666) );
  MXI2XL U1358 ( .A(n5905), .B(n3664), .S0(n369), .Y(n4665) );
  MXI2XL U1359 ( .A(n5904), .B(n3663), .S0(n369), .Y(n4664) );
  MXI2XL U1360 ( .A(n5903), .B(n3662), .S0(n369), .Y(n4663) );
  MXI2XL U1361 ( .A(n5902), .B(n3661), .S0(n369), .Y(n4662) );
  MXI2XL U1362 ( .A(n5901), .B(n3660), .S0(n369), .Y(n4661) );
  MXI2XL U1363 ( .A(n5900), .B(n3659), .S0(n369), .Y(n4660) );
  MXI2XL U1364 ( .A(n5899), .B(n3658), .S0(n369), .Y(n4659) );
  MXI2XL U1365 ( .A(n5898), .B(n3657), .S0(n369), .Y(n4658) );
  MXI2XL U1366 ( .A(n5897), .B(n3656), .S0(n369), .Y(n4657) );
  MXI2XL U1367 ( .A(n5896), .B(n3655), .S0(n369), .Y(n4656) );
  MXI2XL U1368 ( .A(n5895), .B(n3654), .S0(n369), .Y(n4655) );
  MXI2XL U1369 ( .A(n5894), .B(n3653), .S0(n369), .Y(n4654) );
  MXI2XL U1370 ( .A(n5893), .B(n3652), .S0(n369), .Y(n4653) );
  MXI2XL U1371 ( .A(n5892), .B(n3651), .S0(n370), .Y(n4652) );
  MXI2XL U1372 ( .A(n5891), .B(n3650), .S0(n370), .Y(n4651) );
  MXI2XL U1373 ( .A(n5890), .B(n3649), .S0(n370), .Y(n4650) );
  MXI2XL U1374 ( .A(n5889), .B(n3648), .S0(n370), .Y(n4649) );
  MXI2XL U1375 ( .A(n5888), .B(n3647), .S0(n370), .Y(n4648) );
  MXI2XL U1376 ( .A(n5887), .B(n3646), .S0(n370), .Y(n4647) );
  MXI2XL U1377 ( .A(n5886), .B(n3645), .S0(n370), .Y(n4646) );
  MXI2XL U1378 ( .A(n5885), .B(n3644), .S0(n370), .Y(n4645) );
  MXI2XL U1379 ( .A(n5884), .B(n3643), .S0(n370), .Y(n4644) );
  MXI2XL U1380 ( .A(n5883), .B(n3642), .S0(n370), .Y(n4643) );
  MXI2XL U1381 ( .A(n5882), .B(n3641), .S0(n370), .Y(n4642) );
  MXI2XL U1382 ( .A(n5881), .B(n3640), .S0(n370), .Y(n4641) );
  MXI2XL U1383 ( .A(n5880), .B(n3639), .S0(n370), .Y(n4640) );
  MXI2XL U1384 ( .A(n5879), .B(n3638), .S0(n364), .Y(n4639) );
  MXI2XL U1385 ( .A(n5878), .B(n3637), .S0(n366), .Y(n4638) );
  MXI2XL U1386 ( .A(n5877), .B(n3636), .S0(n370), .Y(n4637) );
  MXI2XL U1387 ( .A(n5876), .B(n3635), .S0(n367), .Y(n4636) );
  MXI2XL U1388 ( .A(n5875), .B(n3634), .S0(n371), .Y(n4635) );
  MXI2XL U1389 ( .A(n5751), .B(n3665), .S0(n359), .Y(n4511) );
  MXI2XL U1390 ( .A(n5750), .B(n3664), .S0(n360), .Y(n4510) );
  MXI2XL U1391 ( .A(n5749), .B(n3663), .S0(n360), .Y(n4509) );
  MXI2XL U1392 ( .A(n5748), .B(n3662), .S0(n360), .Y(n4508) );
  MXI2XL U1393 ( .A(n5747), .B(n3661), .S0(n360), .Y(n4507) );
  MXI2XL U1394 ( .A(n5746), .B(n3660), .S0(n360), .Y(n4506) );
  MXI2XL U1395 ( .A(n5745), .B(n3659), .S0(n360), .Y(n4505) );
  MXI2XL U1396 ( .A(n5744), .B(n3658), .S0(n360), .Y(n4504) );
  MXI2XL U1397 ( .A(n5743), .B(n3657), .S0(n360), .Y(n4503) );
  MXI2XL U1398 ( .A(n5742), .B(n3656), .S0(n360), .Y(n4502) );
  MXI2XL U1399 ( .A(n5741), .B(n3655), .S0(n360), .Y(n4501) );
  MXI2XL U1400 ( .A(n5740), .B(n3654), .S0(n360), .Y(n4500) );
  MXI2XL U1401 ( .A(n5739), .B(n3653), .S0(n360), .Y(n4499) );
  MXI2XL U1402 ( .A(n5738), .B(n3652), .S0(n360), .Y(n4498) );
  MXI2XL U1403 ( .A(n5737), .B(n3651), .S0(n361), .Y(n4497) );
  MXI2XL U1404 ( .A(n5736), .B(n3650), .S0(n361), .Y(n4496) );
  MXI2XL U1405 ( .A(n5735), .B(n3649), .S0(n361), .Y(n4495) );
  MXI2XL U1406 ( .A(n5734), .B(n3648), .S0(n361), .Y(n4494) );
  MXI2XL U1407 ( .A(n5733), .B(n3647), .S0(n361), .Y(n4493) );
  MXI2XL U1408 ( .A(n5732), .B(n3646), .S0(n361), .Y(n4492) );
  MXI2XL U1409 ( .A(n5731), .B(n3645), .S0(n361), .Y(n4491) );
  MXI2XL U1410 ( .A(n5730), .B(n3644), .S0(n361), .Y(n4490) );
  MXI2XL U1411 ( .A(n5729), .B(n3643), .S0(n361), .Y(n4489) );
  MXI2XL U1412 ( .A(n5728), .B(n3642), .S0(n361), .Y(n4488) );
  MXI2XL U1413 ( .A(n5727), .B(n3641), .S0(n361), .Y(n4487) );
  MXI2XL U1414 ( .A(n5726), .B(n3640), .S0(n361), .Y(n4486) );
  MXI2XL U1415 ( .A(n5725), .B(n3639), .S0(n361), .Y(n4485) );
  MXI2XL U1416 ( .A(n5724), .B(n3638), .S0(n355), .Y(n4484) );
  MXI2XL U1417 ( .A(n5723), .B(n3637), .S0(n357), .Y(n4483) );
  MXI2XL U1418 ( .A(n5722), .B(n3636), .S0(n361), .Y(n4482) );
  MXI2XL U1419 ( .A(n5721), .B(n3635), .S0(n358), .Y(n4481) );
  MXI2XL U1420 ( .A(n5720), .B(n3634), .S0(n362), .Y(n4480) );
  MXI2XL U1421 ( .A(n5596), .B(n3665), .S0(n349), .Y(n4356) );
  MXI2XL U1422 ( .A(n5595), .B(n3664), .S0(n350), .Y(n4355) );
  MXI2XL U1423 ( .A(n5594), .B(n3663), .S0(n350), .Y(n4354) );
  MXI2XL U1424 ( .A(n5593), .B(n3662), .S0(n350), .Y(n4353) );
  MXI2XL U1425 ( .A(n5592), .B(n3661), .S0(n350), .Y(n4352) );
  MXI2XL U1426 ( .A(n5591), .B(n3660), .S0(n350), .Y(n4351) );
  MXI2XL U1427 ( .A(n5590), .B(n3659), .S0(n350), .Y(n4350) );
  MXI2XL U1428 ( .A(n5589), .B(n3658), .S0(n350), .Y(n4349) );
  MXI2XL U1429 ( .A(n5588), .B(n3657), .S0(n350), .Y(n4348) );
  MXI2XL U1430 ( .A(n5587), .B(n3656), .S0(n350), .Y(n4347) );
  MXI2XL U1431 ( .A(n5586), .B(n3655), .S0(n350), .Y(n4346) );
  MXI2XL U1432 ( .A(n5585), .B(n3654), .S0(n350), .Y(n4345) );
  MXI2XL U1433 ( .A(n5584), .B(n3653), .S0(n350), .Y(n4344) );
  MXI2XL U1434 ( .A(n5583), .B(n3652), .S0(n350), .Y(n4343) );
  MXI2XL U1435 ( .A(n5582), .B(n3651), .S0(n351), .Y(n4342) );
  MXI2XL U1436 ( .A(n5581), .B(n3650), .S0(n351), .Y(n4341) );
  MXI2XL U1437 ( .A(n5580), .B(n3649), .S0(n351), .Y(n4340) );
  MXI2XL U1438 ( .A(n5579), .B(n3648), .S0(n351), .Y(n4339) );
  MXI2XL U1439 ( .A(n5578), .B(n3647), .S0(n351), .Y(n4338) );
  MXI2XL U1440 ( .A(n5577), .B(n3646), .S0(n351), .Y(n4337) );
  MXI2XL U1441 ( .A(n5576), .B(n3645), .S0(n351), .Y(n4336) );
  MXI2XL U1442 ( .A(n5575), .B(n3644), .S0(n351), .Y(n4335) );
  MXI2XL U1443 ( .A(n5574), .B(n3643), .S0(n351), .Y(n4334) );
  MXI2XL U1444 ( .A(n5573), .B(n3642), .S0(n351), .Y(n4333) );
  MXI2XL U1445 ( .A(n5572), .B(n3641), .S0(n351), .Y(n4332) );
  MXI2XL U1446 ( .A(n5571), .B(n3640), .S0(n351), .Y(n4331) );
  MXI2XL U1447 ( .A(n5570), .B(n3639), .S0(n351), .Y(n4330) );
  MXI2XL U1448 ( .A(n5569), .B(n3638), .S0(n345), .Y(n4329) );
  MXI2XL U1449 ( .A(n5568), .B(n3637), .S0(n347), .Y(n4328) );
  MXI2XL U1450 ( .A(n5567), .B(n3636), .S0(n351), .Y(n4327) );
  MXI2XL U1451 ( .A(n5566), .B(n3635), .S0(n348), .Y(n4326) );
  MXI2XL U1452 ( .A(n5565), .B(n3634), .S0(n352), .Y(n4325) );
  MXI2XL U1453 ( .A(n5441), .B(n3665), .S0(n340), .Y(n4201) );
  MXI2XL U1454 ( .A(n5440), .B(n3664), .S0(n341), .Y(n4200) );
  MXI2XL U1455 ( .A(n5439), .B(n3663), .S0(n341), .Y(n4199) );
  MXI2XL U1456 ( .A(n5438), .B(n3662), .S0(n341), .Y(n4198) );
  MXI2XL U1457 ( .A(n5437), .B(n3661), .S0(n341), .Y(n4197) );
  MXI2XL U1458 ( .A(n5436), .B(n3660), .S0(n341), .Y(n4196) );
  MXI2XL U1459 ( .A(n5435), .B(n3659), .S0(n341), .Y(n4195) );
  MXI2XL U1460 ( .A(n5434), .B(n3658), .S0(n341), .Y(n4194) );
  MXI2XL U1461 ( .A(n5433), .B(n3657), .S0(n341), .Y(n4193) );
  MXI2XL U1462 ( .A(n5432), .B(n3656), .S0(n341), .Y(n4192) );
  MXI2XL U1463 ( .A(n5431), .B(n3655), .S0(n341), .Y(n4191) );
  MXI2XL U1464 ( .A(n5430), .B(n3654), .S0(n341), .Y(n4190) );
  MXI2XL U1465 ( .A(n5429), .B(n3653), .S0(n341), .Y(n4189) );
  MXI2XL U1466 ( .A(n5428), .B(n3652), .S0(n341), .Y(n4188) );
  MXI2XL U1467 ( .A(n5427), .B(n3651), .S0(n342), .Y(n4187) );
  MXI2XL U1468 ( .A(n5426), .B(n3650), .S0(n342), .Y(n4186) );
  MXI2XL U1469 ( .A(n5425), .B(n3649), .S0(n342), .Y(n4185) );
  MXI2XL U1470 ( .A(n5424), .B(n3648), .S0(n342), .Y(n4184) );
  MXI2XL U1471 ( .A(n5423), .B(n3647), .S0(n342), .Y(n4183) );
  MXI2XL U1472 ( .A(n5422), .B(n3646), .S0(n342), .Y(n4182) );
  MXI2XL U1473 ( .A(n5421), .B(n3645), .S0(n342), .Y(n4181) );
  MXI2XL U1474 ( .A(n5420), .B(n3644), .S0(n342), .Y(n4180) );
  MXI2XL U1475 ( .A(n5419), .B(n3643), .S0(n342), .Y(n4179) );
  MXI2XL U1476 ( .A(n5418), .B(n3642), .S0(n342), .Y(n4178) );
  MXI2XL U1477 ( .A(n5417), .B(n3641), .S0(n342), .Y(n4177) );
  MXI2XL U1478 ( .A(n5416), .B(n3640), .S0(n342), .Y(n4176) );
  MXI2XL U1479 ( .A(n5415), .B(n3639), .S0(n342), .Y(n4175) );
  MXI2XL U1480 ( .A(n5414), .B(n3638), .S0(n336), .Y(n4174) );
  MXI2XL U1481 ( .A(n5413), .B(n3637), .S0(n338), .Y(n4173) );
  MXI2XL U1482 ( .A(n5412), .B(n3636), .S0(n342), .Y(n4172) );
  MXI2XL U1483 ( .A(n5411), .B(n3635), .S0(n339), .Y(n4171) );
  MXI2XL U1484 ( .A(n5410), .B(n3634), .S0(n343), .Y(n4170) );
  MXI2XL U1485 ( .A(n5286), .B(n3665), .S0(n331), .Y(n4046) );
  MXI2XL U1486 ( .A(n5285), .B(n3664), .S0(n332), .Y(n4045) );
  MXI2XL U1487 ( .A(n5284), .B(n3663), .S0(n332), .Y(n4044) );
  MXI2XL U1488 ( .A(n5283), .B(n3662), .S0(n332), .Y(n4043) );
  MXI2XL U1489 ( .A(n5282), .B(n3661), .S0(n332), .Y(n4042) );
  MXI2XL U1490 ( .A(n5281), .B(n3660), .S0(n332), .Y(n4041) );
  MXI2XL U1491 ( .A(n5280), .B(n3659), .S0(n332), .Y(n4040) );
  MXI2XL U1492 ( .A(n5279), .B(n3658), .S0(n332), .Y(n4039) );
  MXI2XL U1493 ( .A(n5278), .B(n3657), .S0(n332), .Y(n4038) );
  MXI2XL U1494 ( .A(n5277), .B(n3656), .S0(n332), .Y(n4037) );
  MXI2XL U1495 ( .A(n5276), .B(n3655), .S0(n332), .Y(n4036) );
  MXI2XL U1496 ( .A(n5275), .B(n3654), .S0(n332), .Y(n4035) );
  MXI2XL U1497 ( .A(n5274), .B(n3653), .S0(n332), .Y(n4034) );
  MXI2XL U1498 ( .A(n5273), .B(n3652), .S0(n332), .Y(n4033) );
  MXI2XL U1499 ( .A(n5272), .B(n3651), .S0(n333), .Y(n4032) );
  MXI2XL U1500 ( .A(n5271), .B(n3650), .S0(n333), .Y(n4031) );
  MXI2XL U1501 ( .A(n5270), .B(n3649), .S0(n333), .Y(n4030) );
  MXI2XL U1502 ( .A(n5269), .B(n3648), .S0(n333), .Y(n4029) );
  MXI2XL U1503 ( .A(n5268), .B(n3647), .S0(n333), .Y(n4028) );
  MXI2XL U1504 ( .A(n5267), .B(n3646), .S0(n333), .Y(n4027) );
  MXI2XL U1505 ( .A(n5266), .B(n3645), .S0(n333), .Y(n4026) );
  MXI2XL U1506 ( .A(n5265), .B(n3644), .S0(n333), .Y(n4025) );
  MXI2XL U1507 ( .A(n5264), .B(n3643), .S0(n333), .Y(n4024) );
  MXI2XL U1508 ( .A(n5263), .B(n3642), .S0(n333), .Y(n4023) );
  MXI2XL U1509 ( .A(n5262), .B(n3641), .S0(n333), .Y(n4022) );
  MXI2XL U1510 ( .A(n5261), .B(n3640), .S0(n333), .Y(n4021) );
  MXI2XL U1511 ( .A(n5260), .B(n3639), .S0(n333), .Y(n4020) );
  MXI2XL U1512 ( .A(n5259), .B(n3638), .S0(n327), .Y(n4019) );
  MXI2XL U1513 ( .A(n5258), .B(n3637), .S0(n329), .Y(n4018) );
  MXI2XL U1514 ( .A(n5257), .B(n3636), .S0(n333), .Y(n4017) );
  MXI2XL U1515 ( .A(n5256), .B(n3635), .S0(n330), .Y(n4016) );
  MXI2XL U1516 ( .A(n5255), .B(n3634), .S0(n334), .Y(n4015) );
  MXI2XL U1517 ( .A(n5131), .B(n3665), .S0(n322), .Y(n3891) );
  MXI2XL U1518 ( .A(n5130), .B(n3664), .S0(n323), .Y(n3890) );
  MXI2XL U1519 ( .A(n5129), .B(n3663), .S0(n323), .Y(n3889) );
  MXI2XL U1520 ( .A(n5128), .B(n3662), .S0(n323), .Y(n3888) );
  MXI2XL U1521 ( .A(n5127), .B(n3661), .S0(n323), .Y(n3887) );
  MXI2XL U1522 ( .A(n5126), .B(n3660), .S0(n323), .Y(n3886) );
  MXI2XL U1523 ( .A(n5125), .B(n3659), .S0(n323), .Y(n3885) );
  MXI2XL U1524 ( .A(n5124), .B(n3658), .S0(n323), .Y(n3884) );
  MXI2XL U1525 ( .A(n5123), .B(n3657), .S0(n323), .Y(n3883) );
  MXI2XL U1526 ( .A(n5122), .B(n3656), .S0(n323), .Y(n3882) );
  MXI2XL U1527 ( .A(n5121), .B(n3655), .S0(n323), .Y(n3881) );
  MXI2XL U1528 ( .A(n5120), .B(n3654), .S0(n323), .Y(n3880) );
  MXI2XL U1529 ( .A(n5119), .B(n3653), .S0(n323), .Y(n3879) );
  MXI2XL U1530 ( .A(n5118), .B(n3652), .S0(n323), .Y(n3878) );
  MXI2XL U1531 ( .A(n5117), .B(n3651), .S0(n324), .Y(n3877) );
  MXI2XL U1532 ( .A(n5116), .B(n3650), .S0(n324), .Y(n3876) );
  MXI2XL U1533 ( .A(n5115), .B(n3649), .S0(n324), .Y(n3875) );
  MXI2XL U1534 ( .A(n5114), .B(n3648), .S0(n324), .Y(n3874) );
  MXI2XL U1535 ( .A(n5113), .B(n3647), .S0(n324), .Y(n3873) );
  MXI2XL U1536 ( .A(n5112), .B(n3646), .S0(n324), .Y(n3872) );
  MXI2XL U1537 ( .A(n5111), .B(n3645), .S0(n324), .Y(n3871) );
  MXI2XL U1538 ( .A(n5110), .B(n3644), .S0(n324), .Y(n3870) );
  MXI2XL U1539 ( .A(n5109), .B(n3643), .S0(n324), .Y(n3869) );
  MXI2XL U1540 ( .A(n5108), .B(n3642), .S0(n324), .Y(n3868) );
  MXI2XL U1541 ( .A(n5107), .B(n3641), .S0(n324), .Y(n3867) );
  MXI2XL U1542 ( .A(n5106), .B(n3640), .S0(n324), .Y(n3866) );
  MXI2XL U1543 ( .A(n5105), .B(n3639), .S0(n324), .Y(n3865) );
  MXI2XL U1544 ( .A(n5104), .B(n3638), .S0(n318), .Y(n3864) );
  MXI2XL U1545 ( .A(n5103), .B(n3637), .S0(n320), .Y(n3863) );
  MXI2XL U1546 ( .A(n5102), .B(n3636), .S0(n324), .Y(n3862) );
  MXI2XL U1547 ( .A(n5101), .B(n3635), .S0(n321), .Y(n3861) );
  MXI2XL U1548 ( .A(n5100), .B(n3634), .S0(n325), .Y(n3860) );
  MXI2XL U1549 ( .A(n6152), .B(n3601), .S0(n386), .Y(n4912) );
  MXI2XL U1550 ( .A(n6151), .B(n3600), .S0(n390), .Y(n4911) );
  MXI2XL U1551 ( .A(n6150), .B(n3599), .S0(n387), .Y(n4910) );
  MXI2XL U1552 ( .A(n6149), .B(n3598), .S0(n385), .Y(n4909) );
  MXI2XL U1553 ( .A(n6148), .B(n3597), .S0(n389), .Y(n4908) );
  MXI2XL U1554 ( .A(n6147), .B(n3596), .S0(n382), .Y(n4907) );
  MXI2XL U1555 ( .A(n6146), .B(n3595), .S0(n383), .Y(n4906) );
  MXI2XL U1556 ( .A(n6145), .B(n3594), .S0(n386), .Y(n4905) );
  MXI2XL U1557 ( .A(n6144), .B(n3593), .S0(n390), .Y(n4904) );
  MXI2XL U1558 ( .A(n6143), .B(n3592), .S0(n387), .Y(n4903) );
  MXI2XL U1559 ( .A(n6142), .B(n3591), .S0(n385), .Y(n4902) );
  MXI2XL U1560 ( .A(n6141), .B(n3590), .S0(n389), .Y(n4901) );
  MXI2XL U1561 ( .A(n6140), .B(n3589), .S0(n382), .Y(n4900) );
  MXI2XL U1562 ( .A(n6139), .B(n3588), .S0(n383), .Y(n4899) );
  MXI2XL U1563 ( .A(n6138), .B(n3587), .S0(n386), .Y(n4898) );
  MXI2XL U1564 ( .A(n6137), .B(n3586), .S0(n390), .Y(n4897) );
  MXI2XL U1565 ( .A(n6136), .B(n3585), .S0(n390), .Y(n4896) );
  MXI2XL U1566 ( .A(n6135), .B(n3584), .S0(n390), .Y(n4895) );
  MXI2XL U1567 ( .A(n6134), .B(n3583), .S0(n390), .Y(n4894) );
  MXI2XL U1568 ( .A(n6133), .B(n3582), .S0(n390), .Y(n4893) );
  MXI2XL U1569 ( .A(n6132), .B(n3581), .S0(n390), .Y(n4892) );
  MXI2XL U1570 ( .A(n6131), .B(n3580), .S0(n390), .Y(n4891) );
  MXI2XL U1571 ( .A(n6130), .B(n3579), .S0(n390), .Y(n4890) );
  MXI2XL U1572 ( .A(n6129), .B(n3578), .S0(n390), .Y(n4889) );
  MXI2XL U1573 ( .A(n6128), .B(n3577), .S0(n390), .Y(n4888) );
  MXI2XL U1574 ( .A(n5997), .B(n3601), .S0(n377), .Y(n4757) );
  MXI2XL U1575 ( .A(n5996), .B(n3600), .S0(n381), .Y(n4756) );
  MXI2XL U1576 ( .A(n5995), .B(n3599), .S0(n378), .Y(n4755) );
  MXI2XL U1577 ( .A(n5994), .B(n3598), .S0(n376), .Y(n4754) );
  MXI2XL U1578 ( .A(n5993), .B(n3597), .S0(n380), .Y(n4753) );
  MXI2XL U1579 ( .A(n5992), .B(n3596), .S0(n373), .Y(n4752) );
  MXI2XL U1580 ( .A(n5991), .B(n3595), .S0(n374), .Y(n4751) );
  MXI2XL U1581 ( .A(n5990), .B(n3594), .S0(n377), .Y(n4750) );
  MXI2XL U1582 ( .A(n5989), .B(n3593), .S0(n381), .Y(n4749) );
  MXI2XL U1583 ( .A(n5988), .B(n3592), .S0(n378), .Y(n4748) );
  MXI2XL U1584 ( .A(n5987), .B(n3591), .S0(n376), .Y(n4747) );
  MXI2XL U1585 ( .A(n5986), .B(n3590), .S0(n380), .Y(n4746) );
  MXI2XL U1586 ( .A(n5985), .B(n3589), .S0(n373), .Y(n4745) );
  MXI2XL U1587 ( .A(n5984), .B(n3588), .S0(n374), .Y(n4744) );
  MXI2XL U1588 ( .A(n5983), .B(n3587), .S0(n377), .Y(n4743) );
  MXI2XL U1589 ( .A(n5982), .B(n3586), .S0(n381), .Y(n4742) );
  MXI2XL U1590 ( .A(n5981), .B(n3585), .S0(n381), .Y(n4741) );
  MXI2XL U1591 ( .A(n5980), .B(n3584), .S0(n381), .Y(n4740) );
  MXI2XL U1592 ( .A(n5979), .B(n3583), .S0(n381), .Y(n4739) );
  MXI2XL U1593 ( .A(n5978), .B(n3582), .S0(n381), .Y(n4738) );
  MXI2XL U1594 ( .A(n5977), .B(n3581), .S0(n381), .Y(n4737) );
  MXI2XL U1595 ( .A(n5976), .B(n3580), .S0(n381), .Y(n4736) );
  MXI2XL U1596 ( .A(n5975), .B(n3579), .S0(n381), .Y(n4735) );
  MXI2XL U1597 ( .A(n5974), .B(n3578), .S0(n381), .Y(n4734) );
  MXI2XL U1598 ( .A(n5973), .B(n3577), .S0(n381), .Y(n4733) );
  MXI2XL U1599 ( .A(n5842), .B(n3601), .S0(n368), .Y(n4602) );
  MXI2XL U1600 ( .A(n5841), .B(n3600), .S0(n372), .Y(n4601) );
  MXI2XL U1601 ( .A(n5840), .B(n3599), .S0(n369), .Y(n4600) );
  MXI2XL U1602 ( .A(n5839), .B(n3598), .S0(n367), .Y(n4599) );
  MXI2XL U1603 ( .A(n5838), .B(n3597), .S0(n371), .Y(n4598) );
  MXI2XL U1604 ( .A(n5837), .B(n3596), .S0(n364), .Y(n4597) );
  MXI2XL U1605 ( .A(n5836), .B(n3595), .S0(n365), .Y(n4596) );
  MXI2XL U1606 ( .A(n5835), .B(n3594), .S0(n368), .Y(n4595) );
  MXI2XL U1607 ( .A(n5834), .B(n3593), .S0(n372), .Y(n4594) );
  MXI2XL U1608 ( .A(n5833), .B(n3592), .S0(n369), .Y(n4593) );
  MXI2XL U1609 ( .A(n5832), .B(n3591), .S0(n367), .Y(n4592) );
  MXI2XL U1610 ( .A(n5831), .B(n3590), .S0(n371), .Y(n4591) );
  MXI2XL U1611 ( .A(n5830), .B(n3589), .S0(n364), .Y(n4590) );
  MXI2XL U1612 ( .A(n5829), .B(n3588), .S0(n365), .Y(n4589) );
  MXI2XL U1613 ( .A(n5828), .B(n3587), .S0(n368), .Y(n4588) );
  MXI2XL U1614 ( .A(n5827), .B(n3586), .S0(n372), .Y(n4587) );
  MXI2XL U1615 ( .A(n5826), .B(n3585), .S0(n372), .Y(n4586) );
  MXI2XL U1616 ( .A(n5825), .B(n3584), .S0(n372), .Y(n4585) );
  MXI2XL U1617 ( .A(n5824), .B(n3583), .S0(n372), .Y(n4584) );
  MXI2XL U1618 ( .A(n5823), .B(n3582), .S0(n372), .Y(n4583) );
  MXI2XL U1619 ( .A(n5822), .B(n3581), .S0(n372), .Y(n4582) );
  MXI2XL U1620 ( .A(n5821), .B(n3580), .S0(n372), .Y(n4581) );
  MXI2XL U1621 ( .A(n5820), .B(n3579), .S0(n372), .Y(n4580) );
  MXI2XL U1622 ( .A(n5819), .B(n3578), .S0(n372), .Y(n4579) );
  MXI2XL U1623 ( .A(n5818), .B(n3577), .S0(n372), .Y(n4578) );
  MXI2XL U1624 ( .A(n5687), .B(n3601), .S0(n359), .Y(n4447) );
  MXI2XL U1625 ( .A(n5686), .B(n3600), .S0(n363), .Y(n4446) );
  MXI2XL U1626 ( .A(n5685), .B(n3599), .S0(n360), .Y(n4445) );
  MXI2XL U1627 ( .A(n5684), .B(n3598), .S0(n358), .Y(n4444) );
  MXI2XL U1628 ( .A(n5683), .B(n3597), .S0(n362), .Y(n4443) );
  MXI2XL U1629 ( .A(n5682), .B(n3596), .S0(n355), .Y(n4442) );
  MXI2XL U1630 ( .A(n5681), .B(n3595), .S0(n356), .Y(n4441) );
  MXI2XL U1631 ( .A(n5680), .B(n3594), .S0(n359), .Y(n4440) );
  MXI2XL U1632 ( .A(n5679), .B(n3593), .S0(n363), .Y(n4439) );
  MXI2XL U1633 ( .A(n5678), .B(n3592), .S0(n360), .Y(n4438) );
  MXI2XL U1634 ( .A(n5677), .B(n3591), .S0(n358), .Y(n4437) );
  MXI2XL U1635 ( .A(n5676), .B(n3590), .S0(n362), .Y(n4436) );
  MXI2XL U1636 ( .A(n5675), .B(n3589), .S0(n355), .Y(n4435) );
  MXI2XL U1637 ( .A(n5674), .B(n3588), .S0(n356), .Y(n4434) );
  MXI2XL U1638 ( .A(n5673), .B(n3587), .S0(n359), .Y(n4433) );
  MXI2XL U1639 ( .A(n5672), .B(n3586), .S0(n363), .Y(n4432) );
  MXI2XL U1640 ( .A(n5671), .B(n3585), .S0(n363), .Y(n4431) );
  MXI2XL U1641 ( .A(n5670), .B(n3584), .S0(n363), .Y(n4430) );
  MXI2XL U1642 ( .A(n5669), .B(n3583), .S0(n363), .Y(n4429) );
  MXI2XL U1643 ( .A(n5668), .B(n3582), .S0(n363), .Y(n4428) );
  MXI2XL U1644 ( .A(n5667), .B(n3581), .S0(n363), .Y(n4427) );
  MXI2XL U1645 ( .A(n5666), .B(n3580), .S0(n363), .Y(n4426) );
  MXI2XL U1646 ( .A(n5665), .B(n3579), .S0(n363), .Y(n4425) );
  MXI2XL U1647 ( .A(n5664), .B(n3578), .S0(n363), .Y(n4424) );
  MXI2XL U1648 ( .A(n5663), .B(n3577), .S0(n363), .Y(n4423) );
  MXI2XL U1649 ( .A(n5532), .B(n3601), .S0(n349), .Y(n4292) );
  MXI2XL U1650 ( .A(n5531), .B(n3600), .S0(n354), .Y(n4291) );
  MXI2XL U1651 ( .A(n5530), .B(n3599), .S0(n353), .Y(n4290) );
  MXI2XL U1652 ( .A(n5529), .B(n3598), .S0(n353), .Y(n4289) );
  MXI2XL U1653 ( .A(n5528), .B(n3597), .S0(n353), .Y(n4288) );
  MXI2XL U1654 ( .A(n5527), .B(n3596), .S0(n353), .Y(n4287) );
  MXI2XL U1655 ( .A(n5526), .B(n3595), .S0(n353), .Y(n4286) );
  MXI2XL U1656 ( .A(n5525), .B(n3594), .S0(n353), .Y(n4285) );
  MXI2XL U1657 ( .A(n5524), .B(n3593), .S0(n353), .Y(n4284) );
  MXI2XL U1658 ( .A(n5523), .B(n3592), .S0(n353), .Y(n4283) );
  MXI2XL U1659 ( .A(n5522), .B(n3591), .S0(n353), .Y(n4282) );
  MXI2XL U1660 ( .A(n5521), .B(n3590), .S0(n353), .Y(n4281) );
  MXI2XL U1661 ( .A(n5520), .B(n3589), .S0(n353), .Y(n4280) );
  MXI2XL U1662 ( .A(n5519), .B(n3588), .S0(n353), .Y(n4279) );
  MXI2XL U1663 ( .A(n5518), .B(n3587), .S0(n353), .Y(n4278) );
  MXI2XL U1664 ( .A(n5517), .B(n3586), .S0(n354), .Y(n4277) );
  MXI2XL U1665 ( .A(n5516), .B(n3585), .S0(n354), .Y(n4276) );
  MXI2XL U1666 ( .A(n5515), .B(n3584), .S0(n354), .Y(n4275) );
  MXI2XL U1667 ( .A(n5514), .B(n3583), .S0(n354), .Y(n4274) );
  MXI2XL U1668 ( .A(n5513), .B(n3582), .S0(n354), .Y(n4273) );
  MXI2XL U1669 ( .A(n5512), .B(n3581), .S0(n354), .Y(n4272) );
  MXI2XL U1670 ( .A(n5511), .B(n3580), .S0(n354), .Y(n4271) );
  MXI2XL U1671 ( .A(n5510), .B(n3579), .S0(n354), .Y(n4270) );
  MXI2XL U1672 ( .A(n5509), .B(n3578), .S0(n354), .Y(n4269) );
  MXI2XL U1673 ( .A(n5508), .B(n3577), .S0(n354), .Y(n4268) );
  MXI2XL U1674 ( .A(n5377), .B(n3601), .S0(n340), .Y(n4137) );
  MXI2XL U1675 ( .A(n5376), .B(n3600), .S0(n344), .Y(n4136) );
  MXI2XL U1676 ( .A(n5375), .B(n3599), .S0(n341), .Y(n4135) );
  MXI2XL U1677 ( .A(n5374), .B(n3598), .S0(n339), .Y(n4134) );
  MXI2XL U1678 ( .A(n5373), .B(n3597), .S0(n343), .Y(n4133) );
  MXI2XL U1679 ( .A(n5372), .B(n3596), .S0(n336), .Y(n4132) );
  MXI2XL U1680 ( .A(n5371), .B(n3595), .S0(n337), .Y(n4131) );
  MXI2XL U1681 ( .A(n5370), .B(n3594), .S0(n340), .Y(n4130) );
  MXI2XL U1682 ( .A(n5369), .B(n3593), .S0(n344), .Y(n4129) );
  MXI2XL U1683 ( .A(n5368), .B(n3592), .S0(n341), .Y(n4128) );
  MXI2XL U1684 ( .A(n5367), .B(n3591), .S0(n339), .Y(n4127) );
  MXI2XL U1685 ( .A(n5366), .B(n3590), .S0(n343), .Y(n4126) );
  MXI2XL U1686 ( .A(n5365), .B(n3589), .S0(n336), .Y(n4125) );
  MXI2XL U1687 ( .A(n5364), .B(n3588), .S0(n337), .Y(n4124) );
  MXI2XL U1688 ( .A(n5363), .B(n3587), .S0(n340), .Y(n4123) );
  MXI2XL U1689 ( .A(n5362), .B(n3586), .S0(n344), .Y(n4122) );
  MXI2XL U1690 ( .A(n5361), .B(n3585), .S0(n344), .Y(n4121) );
  MXI2XL U1691 ( .A(n5360), .B(n3584), .S0(n344), .Y(n4120) );
  MXI2XL U1692 ( .A(n5359), .B(n3583), .S0(n344), .Y(n4119) );
  MXI2XL U1693 ( .A(n5358), .B(n3582), .S0(n344), .Y(n4118) );
  MXI2XL U1694 ( .A(n5357), .B(n3581), .S0(n344), .Y(n4117) );
  MXI2XL U1695 ( .A(n5356), .B(n3580), .S0(n344), .Y(n4116) );
  MXI2XL U1696 ( .A(n5355), .B(n3579), .S0(n344), .Y(n4115) );
  MXI2XL U1697 ( .A(n5354), .B(n3578), .S0(n344), .Y(n4114) );
  MXI2XL U1698 ( .A(n5353), .B(n3577), .S0(n344), .Y(n4113) );
  MXI2XL U1699 ( .A(n5222), .B(n3601), .S0(n331), .Y(n3982) );
  MXI2XL U1700 ( .A(n5221), .B(n3600), .S0(n335), .Y(n3981) );
  MXI2XL U1701 ( .A(n5220), .B(n3599), .S0(n332), .Y(n3980) );
  MXI2XL U1702 ( .A(n5219), .B(n3598), .S0(n330), .Y(n3979) );
  MXI2XL U1703 ( .A(n5218), .B(n3597), .S0(n334), .Y(n3978) );
  MXI2XL U1704 ( .A(n5217), .B(n3596), .S0(n327), .Y(n3977) );
  MXI2XL U1705 ( .A(n5216), .B(n3595), .S0(n328), .Y(n3976) );
  MXI2XL U1706 ( .A(n5215), .B(n3594), .S0(n331), .Y(n3975) );
  MXI2XL U1707 ( .A(n5214), .B(n3593), .S0(n335), .Y(n3974) );
  MXI2XL U1708 ( .A(n5213), .B(n3592), .S0(n332), .Y(n3973) );
  MXI2XL U1709 ( .A(n5212), .B(n3591), .S0(n330), .Y(n3972) );
  MXI2XL U1710 ( .A(n5211), .B(n3590), .S0(n334), .Y(n3971) );
  MXI2XL U1711 ( .A(n5210), .B(n3589), .S0(n327), .Y(n3970) );
  MXI2XL U1712 ( .A(n5209), .B(n3588), .S0(n328), .Y(n3969) );
  MXI2XL U1713 ( .A(n5208), .B(n3587), .S0(n331), .Y(n3968) );
  MXI2XL U1714 ( .A(n5207), .B(n3586), .S0(n335), .Y(n3967) );
  MXI2XL U1715 ( .A(n5206), .B(n3585), .S0(n335), .Y(n3966) );
  MXI2XL U1716 ( .A(n5205), .B(n3584), .S0(n335), .Y(n3965) );
  MXI2XL U1717 ( .A(n5204), .B(n3583), .S0(n335), .Y(n3964) );
  MXI2XL U1718 ( .A(n5203), .B(n3582), .S0(n335), .Y(n3963) );
  MXI2XL U1719 ( .A(n5202), .B(n3581), .S0(n335), .Y(n3962) );
  MXI2XL U1720 ( .A(n5201), .B(n3580), .S0(n335), .Y(n3961) );
  MXI2XL U1721 ( .A(n5200), .B(n3579), .S0(n335), .Y(n3960) );
  MXI2XL U1722 ( .A(n5199), .B(n3578), .S0(n335), .Y(n3959) );
  MXI2XL U1723 ( .A(n5198), .B(n3577), .S0(n335), .Y(n3958) );
  MXI2XL U1724 ( .A(n5067), .B(n3601), .S0(n322), .Y(n3827) );
  MXI2XL U1725 ( .A(n5066), .B(n3600), .S0(n326), .Y(n3826) );
  MXI2XL U1726 ( .A(n5065), .B(n3599), .S0(n323), .Y(n3825) );
  MXI2XL U1727 ( .A(n5064), .B(n3598), .S0(n321), .Y(n3824) );
  MXI2XL U1728 ( .A(n5063), .B(n3597), .S0(n325), .Y(n3823) );
  MXI2XL U1729 ( .A(n5062), .B(n3596), .S0(n318), .Y(n3822) );
  MXI2XL U1730 ( .A(n5061), .B(n3595), .S0(n319), .Y(n3821) );
  MXI2XL U1731 ( .A(n5060), .B(n3594), .S0(n322), .Y(n3820) );
  MXI2XL U1732 ( .A(n5059), .B(n3593), .S0(n326), .Y(n3819) );
  MXI2XL U1733 ( .A(n5058), .B(n3592), .S0(n323), .Y(n3818) );
  MXI2XL U1734 ( .A(n5057), .B(n3591), .S0(n321), .Y(n3817) );
  MXI2XL U1735 ( .A(n5056), .B(n3590), .S0(n325), .Y(n3816) );
  MXI2XL U1736 ( .A(n5055), .B(n3589), .S0(n318), .Y(n3815) );
  MXI2XL U1737 ( .A(n5054), .B(n3588), .S0(n319), .Y(n3814) );
  MXI2XL U1738 ( .A(n5053), .B(n3587), .S0(n322), .Y(n3813) );
  MXI2XL U1739 ( .A(n5052), .B(n3586), .S0(n326), .Y(n3812) );
  MXI2XL U1740 ( .A(n5051), .B(n3585), .S0(n326), .Y(n3811) );
  MXI2XL U1741 ( .A(n5050), .B(n3584), .S0(n326), .Y(n3810) );
  MXI2XL U1742 ( .A(n5049), .B(n3583), .S0(n326), .Y(n3809) );
  MXI2XL U1743 ( .A(n5048), .B(n3582), .S0(n326), .Y(n3808) );
  MXI2XL U1744 ( .A(n5047), .B(n3581), .S0(n326), .Y(n3807) );
  MXI2XL U1745 ( .A(n5046), .B(n3580), .S0(n326), .Y(n3806) );
  MXI2XL U1746 ( .A(n5045), .B(n3579), .S0(n326), .Y(n3805) );
  MXI2XL U1747 ( .A(n5044), .B(n3578), .S0(n326), .Y(n3804) );
  MXI2XL U1748 ( .A(n5043), .B(n3577), .S0(n326), .Y(n3803) );
  MXI2XL U1749 ( .A(n6126), .B(n3574), .S0(n390), .Y(n4886) );
  MXI2XL U1750 ( .A(n5971), .B(n3574), .S0(n381), .Y(n4731) );
  MXI2XL U1751 ( .A(n5816), .B(n3574), .S0(n372), .Y(n4576) );
  MXI2XL U1752 ( .A(n5661), .B(n3574), .S0(n363), .Y(n4421) );
  MXI2XL U1753 ( .A(n5506), .B(n3574), .S0(n354), .Y(n4266) );
  MXI2XL U1754 ( .A(n5351), .B(n3574), .S0(n344), .Y(n4111) );
  MXI2XL U1755 ( .A(n5196), .B(n3574), .S0(n335), .Y(n3956) );
  MXI2XL U1756 ( .A(n5041), .B(n3574), .S0(n326), .Y(n3801) );
  MXI2XL U1757 ( .A(n6127), .B(n3576), .S0(n390), .Y(n4887) );
  MXI2XL U1758 ( .A(n5972), .B(n3576), .S0(n381), .Y(n4732) );
  MXI2XL U1759 ( .A(n5817), .B(n3576), .S0(n372), .Y(n4577) );
  MXI2XL U1760 ( .A(n5662), .B(n3576), .S0(n363), .Y(n4422) );
  MXI2XL U1761 ( .A(n5507), .B(n3576), .S0(n354), .Y(n4267) );
  MXI2XL U1762 ( .A(n5352), .B(n3576), .S0(n344), .Y(n4112) );
  MXI2XL U1763 ( .A(n5197), .B(n3576), .S0(n335), .Y(n3957) );
  MXI2XL U1764 ( .A(n5042), .B(n3576), .S0(n326), .Y(n3802) );
  CLKINVX1 U1765 ( .A(proc_reset), .Y(n3094) );
  CLKINVX1 U1766 ( .A(N31), .Y(n461) );
  CLKINVX1 U1767 ( .A(N30), .Y(n437) );
  CLKINVX1 U1768 ( .A(N32), .Y(n473) );
  CLKBUFX3 U1769 ( .A(n390), .Y(n382) );
  CLKBUFX3 U1770 ( .A(n390), .Y(n383) );
  CLKBUFX3 U1771 ( .A(n390), .Y(n384) );
  CLKBUFX3 U1772 ( .A(n387), .Y(n385) );
  CLKBUFX3 U1773 ( .A(n390), .Y(n386) );
  CLKBUFX3 U1774 ( .A(n3736), .Y(n387) );
  CLKBUFX3 U1775 ( .A(n387), .Y(n388) );
  CLKBUFX3 U1776 ( .A(n387), .Y(n389) );
  CLKBUFX3 U1777 ( .A(n381), .Y(n373) );
  CLKBUFX3 U1778 ( .A(n381), .Y(n374) );
  CLKBUFX3 U1779 ( .A(n381), .Y(n375) );
  CLKBUFX3 U1780 ( .A(n378), .Y(n376) );
  CLKBUFX3 U1781 ( .A(n381), .Y(n377) );
  CLKBUFX3 U1782 ( .A(n3735), .Y(n378) );
  CLKBUFX3 U1783 ( .A(n378), .Y(n379) );
  CLKBUFX3 U1784 ( .A(n378), .Y(n380) );
  CLKBUFX3 U1785 ( .A(n372), .Y(n364) );
  CLKBUFX3 U1786 ( .A(n372), .Y(n365) );
  CLKBUFX3 U1787 ( .A(n372), .Y(n366) );
  CLKBUFX3 U1788 ( .A(n369), .Y(n367) );
  CLKBUFX3 U1789 ( .A(n372), .Y(n368) );
  CLKBUFX3 U1790 ( .A(n3734), .Y(n369) );
  CLKBUFX3 U1791 ( .A(n369), .Y(n370) );
  CLKBUFX3 U1792 ( .A(n369), .Y(n371) );
  CLKBUFX3 U1793 ( .A(n363), .Y(n355) );
  CLKBUFX3 U1794 ( .A(n363), .Y(n356) );
  CLKBUFX3 U1795 ( .A(n363), .Y(n357) );
  CLKBUFX3 U1796 ( .A(n360), .Y(n358) );
  CLKBUFX3 U1797 ( .A(n363), .Y(n359) );
  CLKBUFX3 U1798 ( .A(n3733), .Y(n360) );
  CLKBUFX3 U1799 ( .A(n360), .Y(n361) );
  CLKBUFX3 U1800 ( .A(n360), .Y(n362) );
  CLKBUFX3 U1801 ( .A(n3736), .Y(n390) );
  CLKBUFX3 U1802 ( .A(n3735), .Y(n381) );
  CLKBUFX3 U1803 ( .A(n3734), .Y(n372) );
  CLKBUFX3 U1804 ( .A(n3733), .Y(n363) );
  CLKBUFX3 U1805 ( .A(n3058), .Y(n3055) );
  CLKBUFX3 U1806 ( .A(n3058), .Y(n3056) );
  CLKBUFX3 U1807 ( .A(n3074), .Y(n511) );
  CLKBUFX3 U1808 ( .A(n3074), .Y(n510) );
  CLKBUFX3 U1809 ( .A(n3075), .Y(n509) );
  CLKBUFX3 U1810 ( .A(n3075), .Y(n508) );
  CLKBUFX3 U1811 ( .A(n3075), .Y(n507) );
  CLKBUFX3 U1812 ( .A(n3075), .Y(n506) );
  CLKBUFX3 U1813 ( .A(n3076), .Y(n505) );
  CLKBUFX3 U1814 ( .A(n3076), .Y(n504) );
  CLKBUFX3 U1815 ( .A(n3076), .Y(n503) );
  CLKBUFX3 U1816 ( .A(n3076), .Y(n502) );
  CLKBUFX3 U1817 ( .A(n3077), .Y(n501) );
  CLKBUFX3 U1818 ( .A(n3077), .Y(n500) );
  CLKBUFX3 U1819 ( .A(n3077), .Y(n499) );
  CLKBUFX3 U1820 ( .A(n3077), .Y(n498) );
  CLKBUFX3 U1821 ( .A(n3078), .Y(n497) );
  CLKBUFX3 U1822 ( .A(n3078), .Y(n496) );
  CLKBUFX3 U1823 ( .A(n3078), .Y(n495) );
  CLKBUFX3 U1824 ( .A(n3078), .Y(n494) );
  CLKBUFX3 U1825 ( .A(n3079), .Y(n493) );
  CLKBUFX3 U1826 ( .A(n3079), .Y(n492) );
  CLKBUFX3 U1827 ( .A(n3069), .Y(n532) );
  CLKBUFX3 U1828 ( .A(n3069), .Y(n531) );
  CLKBUFX3 U1829 ( .A(n3069), .Y(n530) );
  CLKBUFX3 U1830 ( .A(n3070), .Y(n529) );
  CLKBUFX3 U1831 ( .A(n3070), .Y(n528) );
  CLKBUFX3 U1832 ( .A(n3070), .Y(n527) );
  CLKBUFX3 U1833 ( .A(n3070), .Y(n526) );
  CLKBUFX3 U1834 ( .A(n3071), .Y(n525) );
  CLKBUFX3 U1835 ( .A(n3071), .Y(n524) );
  CLKBUFX3 U1836 ( .A(n3071), .Y(n523) );
  CLKBUFX3 U1837 ( .A(n3071), .Y(n522) );
  CLKBUFX3 U1838 ( .A(n3072), .Y(n521) );
  CLKBUFX3 U1839 ( .A(n3072), .Y(n520) );
  CLKBUFX3 U1840 ( .A(n3072), .Y(n519) );
  CLKBUFX3 U1841 ( .A(n3072), .Y(n518) );
  CLKBUFX3 U1842 ( .A(n3073), .Y(n517) );
  CLKBUFX3 U1843 ( .A(n3073), .Y(n516) );
  CLKBUFX3 U1844 ( .A(n3073), .Y(n515) );
  CLKBUFX3 U1845 ( .A(n3073), .Y(n514) );
  CLKBUFX3 U1846 ( .A(n3074), .Y(n513) );
  CLKBUFX3 U1847 ( .A(n3074), .Y(n512) );
  CLKBUFX3 U1848 ( .A(n3058), .Y(n3054) );
  CLKBUFX3 U1849 ( .A(n3059), .Y(n3053) );
  CLKBUFX3 U1850 ( .A(n3059), .Y(n3052) );
  CLKBUFX3 U1851 ( .A(n3059), .Y(n3051) );
  CLKBUFX3 U1852 ( .A(n3059), .Y(n3050) );
  CLKBUFX3 U1853 ( .A(n3060), .Y(n3049) );
  CLKBUFX3 U1854 ( .A(n3060), .Y(n3048) );
  CLKBUFX3 U1855 ( .A(n3060), .Y(n3047) );
  CLKBUFX3 U1856 ( .A(n3060), .Y(n3046) );
  CLKBUFX3 U1857 ( .A(n3061), .Y(n3045) );
  CLKBUFX3 U1858 ( .A(n3061), .Y(n3044) );
  CLKBUFX3 U1859 ( .A(n3061), .Y(n3043) );
  CLKBUFX3 U1860 ( .A(n3061), .Y(n3042) );
  CLKBUFX3 U1861 ( .A(n3062), .Y(n3041) );
  CLKBUFX3 U1862 ( .A(n3062), .Y(n3040) );
  CLKBUFX3 U1863 ( .A(n3062), .Y(n3039) );
  CLKBUFX3 U1864 ( .A(n3062), .Y(n3038) );
  CLKBUFX3 U1865 ( .A(n3063), .Y(n3037) );
  CLKBUFX3 U1866 ( .A(n3063), .Y(n3036) );
  CLKBUFX3 U1867 ( .A(n3063), .Y(n3035) );
  CLKBUFX3 U1868 ( .A(n3063), .Y(n3034) );
  CLKBUFX3 U1869 ( .A(n3064), .Y(n3033) );
  CLKBUFX3 U1870 ( .A(n3064), .Y(n3032) );
  CLKBUFX3 U1871 ( .A(n3064), .Y(n3031) );
  CLKBUFX3 U1872 ( .A(n3064), .Y(n3030) );
  CLKBUFX3 U1873 ( .A(n3065), .Y(n3029) );
  CLKBUFX3 U1874 ( .A(n3065), .Y(n3028) );
  CLKBUFX3 U1875 ( .A(n3065), .Y(n3027) );
  CLKBUFX3 U1876 ( .A(n3065), .Y(n3026) );
  CLKBUFX3 U1877 ( .A(n3066), .Y(n3025) );
  CLKBUFX3 U1878 ( .A(n3066), .Y(n3024) );
  CLKBUFX3 U1879 ( .A(n3066), .Y(n3023) );
  CLKBUFX3 U1880 ( .A(n3066), .Y(n3022) );
  CLKBUFX3 U1881 ( .A(n3067), .Y(n3020) );
  CLKBUFX3 U1882 ( .A(n3067), .Y(n540) );
  CLKBUFX3 U1883 ( .A(n3067), .Y(n539) );
  CLKBUFX3 U1884 ( .A(n3067), .Y(n538) );
  CLKBUFX3 U1885 ( .A(n3068), .Y(n537) );
  CLKBUFX3 U1886 ( .A(n3068), .Y(n536) );
  CLKBUFX3 U1887 ( .A(n3068), .Y(n535) );
  CLKBUFX3 U1888 ( .A(n3068), .Y(n534) );
  CLKBUFX3 U1889 ( .A(n3069), .Y(n533) );
  CLKBUFX3 U1890 ( .A(n3079), .Y(n491) );
  CLKBUFX3 U1891 ( .A(n3080), .Y(n489) );
  CLKBUFX3 U1892 ( .A(n3080), .Y(n488) );
  CLKBUFX3 U1893 ( .A(n3080), .Y(n487) );
  CLKBUFX3 U1894 ( .A(n3080), .Y(n486) );
  CLKBUFX3 U1895 ( .A(n3081), .Y(n485) );
  CLKBUFX3 U1896 ( .A(n3081), .Y(n484) );
  CLKBUFX3 U1897 ( .A(n3081), .Y(n483) );
  CLKBUFX3 U1898 ( .A(n3079), .Y(n490) );
  CLKBUFX3 U1899 ( .A(n3081), .Y(n482) );
  CLKBUFX3 U1900 ( .A(n354), .Y(n345) );
  CLKBUFX3 U1901 ( .A(n354), .Y(n346) );
  CLKBUFX3 U1902 ( .A(n353), .Y(n347) );
  CLKBUFX3 U1903 ( .A(n350), .Y(n348) );
  CLKBUFX3 U1904 ( .A(n354), .Y(n349) );
  CLKBUFX3 U1905 ( .A(n3732), .Y(n350) );
  CLKBUFX3 U1906 ( .A(n353), .Y(n351) );
  CLKBUFX3 U1907 ( .A(n350), .Y(n352) );
  CLKBUFX3 U1908 ( .A(n3732), .Y(n353) );
  CLKBUFX3 U1909 ( .A(n344), .Y(n336) );
  CLKBUFX3 U1910 ( .A(n344), .Y(n337) );
  CLKBUFX3 U1911 ( .A(n344), .Y(n338) );
  CLKBUFX3 U1912 ( .A(n341), .Y(n339) );
  CLKBUFX3 U1913 ( .A(n344), .Y(n340) );
  CLKBUFX3 U1914 ( .A(n3731), .Y(n341) );
  CLKBUFX3 U1915 ( .A(n341), .Y(n342) );
  CLKBUFX3 U1916 ( .A(n341), .Y(n343) );
  CLKBUFX3 U1917 ( .A(n335), .Y(n327) );
  CLKBUFX3 U1918 ( .A(n335), .Y(n328) );
  CLKBUFX3 U1919 ( .A(n335), .Y(n329) );
  CLKBUFX3 U1920 ( .A(n332), .Y(n330) );
  CLKBUFX3 U1921 ( .A(n335), .Y(n331) );
  CLKBUFX3 U1922 ( .A(n3730), .Y(n332) );
  CLKBUFX3 U1923 ( .A(n332), .Y(n333) );
  CLKBUFX3 U1924 ( .A(n332), .Y(n334) );
  CLKBUFX3 U1925 ( .A(n326), .Y(n318) );
  CLKBUFX3 U1926 ( .A(n326), .Y(n319) );
  CLKBUFX3 U1927 ( .A(n326), .Y(n320) );
  CLKBUFX3 U1928 ( .A(n323), .Y(n321) );
  CLKBUFX3 U1929 ( .A(n326), .Y(n322) );
  CLKBUFX3 U1930 ( .A(n3575), .Y(n323) );
  CLKBUFX3 U1931 ( .A(n323), .Y(n324) );
  CLKBUFX3 U1932 ( .A(n323), .Y(n325) );
  CLKBUFX3 U1933 ( .A(n3732), .Y(n354) );
  CLKBUFX3 U1934 ( .A(n3731), .Y(n344) );
  CLKBUFX3 U1935 ( .A(n3730), .Y(n335) );
  CLKBUFX3 U1936 ( .A(n3575), .Y(n326) );
  INVX3 U1937 ( .A(n413), .Y(n402) );
  INVX3 U1938 ( .A(n413), .Y(n403) );
  INVX3 U1939 ( .A(n413), .Y(n404) );
  INVX3 U1940 ( .A(n413), .Y(n405) );
  INVX3 U1941 ( .A(n414), .Y(n406) );
  INVX3 U1942 ( .A(n315), .Y(n407) );
  INVX3 U1943 ( .A(n410), .Y(n399) );
  INVX3 U1944 ( .A(n413), .Y(n400) );
  INVX3 U1945 ( .A(n315), .Y(n401) );
  INVX3 U1946 ( .A(n410), .Y(n408) );
  CLKBUFX3 U1947 ( .A(n3058), .Y(n3057) );
  INVX3 U1948 ( .A(n414), .Y(n409) );
  CLKBUFX3 U1949 ( .A(n3082), .Y(n481) );
  CLKBUFX3 U1950 ( .A(n3082), .Y(n480) );
  CLKBUFX3 U1951 ( .A(n3082), .Y(n479) );
  CLKBUFX3 U1952 ( .A(n3082), .Y(n478) );
  CLKBUFX3 U1953 ( .A(n3083), .Y(n477) );
  CLKBUFX3 U1954 ( .A(n3083), .Y(n476) );
  CLKBUFX3 U1955 ( .A(n3083), .Y(n475) );
  CLKBUFX3 U1956 ( .A(n3083), .Y(n474) );
  CLKBUFX3 U1957 ( .A(n414), .Y(n412) );
  CLKBUFX3 U1958 ( .A(n315), .Y(n410) );
  CLKBUFX3 U1959 ( .A(n414), .Y(mem_write) );
  CLKBUFX3 U1960 ( .A(n3092), .Y(n3075) );
  CLKBUFX3 U1961 ( .A(n3085), .Y(n3076) );
  CLKBUFX3 U1962 ( .A(n3085), .Y(n3077) );
  CLKBUFX3 U1963 ( .A(n3084), .Y(n3078) );
  CLKBUFX3 U1964 ( .A(n3086), .Y(n3070) );
  CLKBUFX3 U1965 ( .A(n3086), .Y(n3071) );
  CLKBUFX3 U1966 ( .A(n3091), .Y(n3072) );
  CLKBUFX3 U1967 ( .A(n3091), .Y(n3073) );
  CLKBUFX3 U1968 ( .A(n3092), .Y(n3074) );
  CLKBUFX3 U1969 ( .A(n3088), .Y(n3059) );
  CLKBUFX3 U1970 ( .A(n3088), .Y(n3060) );
  CLKBUFX3 U1971 ( .A(n3087), .Y(n3061) );
  CLKBUFX3 U1972 ( .A(n3089), .Y(n3062) );
  CLKBUFX3 U1973 ( .A(n3085), .Y(n3063) );
  CLKBUFX3 U1974 ( .A(n3089), .Y(n3064) );
  CLKBUFX3 U1975 ( .A(n3086), .Y(n3065) );
  CLKBUFX3 U1976 ( .A(n3087), .Y(n3066) );
  CLKBUFX3 U1977 ( .A(n3087), .Y(n3067) );
  CLKBUFX3 U1978 ( .A(n3090), .Y(n3068) );
  CLKBUFX3 U1979 ( .A(n3090), .Y(n3069) );
  CLKBUFX3 U1980 ( .A(n3093), .Y(n3080) );
  CLKBUFX3 U1981 ( .A(n3084), .Y(n3079) );
  CLKBUFX3 U1982 ( .A(n3093), .Y(n3081) );
  CLKBUFX3 U1983 ( .A(n3088), .Y(n3058) );
  INVX3 U1984 ( .A(n436), .Y(n423) );
  INVX3 U1985 ( .A(n436), .Y(n417) );
  INVX3 U1986 ( .A(n435), .Y(n424) );
  INVX3 U1987 ( .A(n435), .Y(n418) );
  INVX3 U1988 ( .A(n435), .Y(n425) );
  INVX3 U1989 ( .A(n436), .Y(n426) );
  INVX3 U1990 ( .A(n436), .Y(n427) );
  INVX3 U1991 ( .A(n435), .Y(n428) );
  INVX3 U1992 ( .A(n435), .Y(n429) );
  INVX3 U1993 ( .A(n437), .Y(n430) );
  INVX3 U1994 ( .A(n437), .Y(n431) );
  INVX3 U1995 ( .A(n435), .Y(n432) );
  INVX3 U1996 ( .A(n435), .Y(n433) );
  INVX3 U1997 ( .A(n435), .Y(n415) );
  INVX3 U1998 ( .A(n435), .Y(n416) );
  INVX3 U1999 ( .A(n435), .Y(n419) );
  INVX3 U2000 ( .A(n436), .Y(n420) );
  INVX3 U2001 ( .A(n436), .Y(n421) );
  INVX3 U2002 ( .A(n436), .Y(n422) );
  INVX3 U2003 ( .A(n459), .Y(n458) );
  INVX3 U2004 ( .A(n460), .Y(n438) );
  INVX3 U2005 ( .A(n459), .Y(n439) );
  INVX3 U2006 ( .A(n460), .Y(n440) );
  INVX3 U2007 ( .A(n459), .Y(n441) );
  INVX3 U2008 ( .A(n459), .Y(n442) );
  INVX3 U2009 ( .A(n460), .Y(n443) );
  INVX3 U2010 ( .A(n459), .Y(n444) );
  INVX3 U2011 ( .A(n460), .Y(n445) );
  INVX3 U2012 ( .A(n460), .Y(n446) );
  INVX3 U2013 ( .A(n460), .Y(n447) );
  INVX3 U2014 ( .A(n460), .Y(n448) );
  INVX3 U2015 ( .A(n460), .Y(n451) );
  INVX3 U2016 ( .A(n461), .Y(n452) );
  INVX3 U2017 ( .A(n459), .Y(n453) );
  INVX3 U2018 ( .A(n460), .Y(n454) );
  INVX3 U2019 ( .A(n460), .Y(n449) );
  INVX3 U2020 ( .A(n461), .Y(n450) );
  INVX3 U2021 ( .A(n459), .Y(n455) );
  INVX3 U2022 ( .A(n459), .Y(n456) );
  INVX3 U2023 ( .A(n459), .Y(n457) );
  CLKBUFX3 U2024 ( .A(n395), .Y(n396) );
  CLKBUFX3 U2025 ( .A(n3741), .Y(n395) );
  CLKBUFX3 U2026 ( .A(n3741), .Y(n394) );
  CLKBUFX3 U2027 ( .A(n3741), .Y(n393) );
  CLKBUFX3 U2028 ( .A(n393), .Y(n397) );
  CLKBUFX3 U2029 ( .A(n3741), .Y(n398) );
  CLKBUFX3 U2030 ( .A(n395), .Y(n392) );
  CLKBUFX3 U2031 ( .A(n414), .Y(n413) );
  CLKBUFX3 U2032 ( .A(n3092), .Y(n3085) );
  CLKBUFX3 U2033 ( .A(n3091), .Y(n3086) );
  CLKBUFX3 U2034 ( .A(n3090), .Y(n3087) );
  CLKBUFX3 U2035 ( .A(n3093), .Y(n3084) );
  CLKBUFX3 U2036 ( .A(n3095), .Y(n3082) );
  CLKBUFX3 U2037 ( .A(n3089), .Y(n3083) );
  INVX3 U2038 ( .A(n436), .Y(n434) );
  INVX3 U2039 ( .A(n473), .Y(n470) );
  INVX3 U2040 ( .A(n472), .Y(n462) );
  INVX3 U2041 ( .A(n472), .Y(n466) );
  INVX3 U2042 ( .A(n472), .Y(n463) );
  INVX3 U2043 ( .A(n472), .Y(n467) );
  INVX3 U2044 ( .A(n472), .Y(n464) );
  INVX3 U2045 ( .A(n473), .Y(n465) );
  INVX3 U2046 ( .A(n472), .Y(n468) );
  INVX3 U2047 ( .A(n473), .Y(n469) );
  CLKBUFX3 U2048 ( .A(n437), .Y(n435) );
  CLKBUFX3 U2049 ( .A(n460), .Y(n459) );
  CLKBUFX3 U2050 ( .A(n437), .Y(n436) );
  CLKBUFX3 U2051 ( .A(n461), .Y(n460) );
  CLKBUFX3 U2052 ( .A(n3094), .Y(n3091) );
  CLKBUFX3 U2053 ( .A(n3094), .Y(n3092) );
  CLKBUFX3 U2054 ( .A(n3094), .Y(n3090) );
  CLKBUFX3 U2055 ( .A(n3094), .Y(n3093) );
  CLKBUFX3 U2056 ( .A(n3095), .Y(n3089) );
  CLKBUFX3 U2057 ( .A(n3095), .Y(n3088) );
  CLKBUFX3 U2058 ( .A(n315), .Y(n414) );
  CLKINVX1 U2059 ( .A(n472), .Y(n471) );
  INVX1 U2060 ( .A(proc_reset), .Y(n3095) );
  AND4X1 U2061 ( .A(N34), .B(n3767), .C(n3760), .D(n3740), .Y(n315) );
  CLKBUFX3 U2062 ( .A(n473), .Y(n472) );
  CLKMX2X2 U2063 ( .A(n316), .B(n317), .S0(n470), .Y(N34) );
  MX4X1 U2064 ( .A(\CACHE[0][153] ), .B(\CACHE[1][153] ), .C(\CACHE[2][153] ), 
        .D(\CACHE[3][153] ), .S0(n421), .S1(n458), .Y(n316) );
  MX4X1 U2065 ( .A(\CACHE[4][153] ), .B(\CACHE[5][153] ), .C(\CACHE[6][153] ), 
        .D(\CACHE[7][153] ), .S0(n434), .S1(n458), .Y(n317) );
  MXI2X1 U2066 ( .A(n3358), .B(n3359), .S0(n468), .Y(N56) );
  MXI4X1 U2067 ( .A(\CACHE[4][131] ), .B(\CACHE[5][131] ), .C(\CACHE[6][131] ), 
        .D(\CACHE[7][131] ), .S0(n420), .S1(n455), .Y(n3359) );
  MXI4X1 U2068 ( .A(\CACHE[0][131] ), .B(\CACHE[1][131] ), .C(\CACHE[2][131] ), 
        .D(\CACHE[3][131] ), .S0(n420), .S1(n455), .Y(n3358) );
  MXI2X1 U2069 ( .A(n3360), .B(n3361), .S0(n469), .Y(N55) );
  MXI4X1 U2070 ( .A(\CACHE[4][132] ), .B(\CACHE[5][132] ), .C(\CACHE[6][132] ), 
        .D(\CACHE[7][132] ), .S0(n420), .S1(n440), .Y(n3361) );
  MXI4X1 U2071 ( .A(\CACHE[0][132] ), .B(\CACHE[1][132] ), .C(\CACHE[2][132] ), 
        .D(\CACHE[3][132] ), .S0(n420), .S1(n438), .Y(n3360) );
  MXI2X1 U2072 ( .A(n3362), .B(n3363), .S0(n469), .Y(N54) );
  MXI4X1 U2073 ( .A(\CACHE[4][133] ), .B(\CACHE[5][133] ), .C(\CACHE[6][133] ), 
        .D(\CACHE[7][133] ), .S0(n420), .S1(n451), .Y(n3363) );
  MXI4X1 U2074 ( .A(\CACHE[0][133] ), .B(\CACHE[1][133] ), .C(\CACHE[2][133] ), 
        .D(\CACHE[3][133] ), .S0(n420), .S1(n448), .Y(n3362) );
  MXI2X1 U2075 ( .A(n3370), .B(n3371), .S0(n469), .Y(N50) );
  MXI4X1 U2076 ( .A(\CACHE[4][137] ), .B(\CACHE[5][137] ), .C(\CACHE[6][137] ), 
        .D(\CACHE[7][137] ), .S0(n421), .S1(n439), .Y(n3371) );
  MXI4X1 U2077 ( .A(\CACHE[0][137] ), .B(\CACHE[1][137] ), .C(\CACHE[2][137] ), 
        .D(\CACHE[3][137] ), .S0(n421), .S1(n456), .Y(n3370) );
  MXI2X1 U2078 ( .A(n3372), .B(n3373), .S0(n469), .Y(N49) );
  MXI4X1 U2079 ( .A(\CACHE[4][138] ), .B(\CACHE[5][138] ), .C(\CACHE[6][138] ), 
        .D(\CACHE[7][138] ), .S0(n421), .S1(n456), .Y(n3373) );
  MXI4X1 U2080 ( .A(\CACHE[0][138] ), .B(\CACHE[1][138] ), .C(\CACHE[2][138] ), 
        .D(\CACHE[3][138] ), .S0(n421), .S1(n456), .Y(n3372) );
  MXI2X1 U2081 ( .A(n3374), .B(n3375), .S0(n469), .Y(N48) );
  MXI4X1 U2082 ( .A(\CACHE[4][139] ), .B(\CACHE[5][139] ), .C(\CACHE[6][139] ), 
        .D(\CACHE[7][139] ), .S0(n421), .S1(n456), .Y(n3375) );
  MXI4X1 U2083 ( .A(\CACHE[0][139] ), .B(\CACHE[1][139] ), .C(\CACHE[2][139] ), 
        .D(\CACHE[3][139] ), .S0(n421), .S1(n456), .Y(n3374) );
  MXI2X1 U2084 ( .A(n3382), .B(n3383), .S0(n469), .Y(N44) );
  MXI4X1 U2085 ( .A(\CACHE[4][143] ), .B(\CACHE[5][143] ), .C(\CACHE[6][143] ), 
        .D(\CACHE[7][143] ), .S0(n422), .S1(n456), .Y(n3383) );
  MXI4X1 U2086 ( .A(\CACHE[0][143] ), .B(\CACHE[1][143] ), .C(\CACHE[2][143] ), 
        .D(\CACHE[3][143] ), .S0(n422), .S1(n456), .Y(n3382) );
  MXI2X1 U2087 ( .A(n3384), .B(n3385), .S0(n470), .Y(N43) );
  MXI4X1 U2088 ( .A(\CACHE[4][144] ), .B(\CACHE[5][144] ), .C(\CACHE[6][144] ), 
        .D(\CACHE[7][144] ), .S0(n422), .S1(n457), .Y(n3385) );
  MXI4X1 U2089 ( .A(\CACHE[0][144] ), .B(\CACHE[1][144] ), .C(\CACHE[2][144] ), 
        .D(\CACHE[3][144] ), .S0(n422), .S1(n457), .Y(n3384) );
  MXI2X1 U2090 ( .A(n3386), .B(n3387), .S0(n470), .Y(N42) );
  MXI4X1 U2091 ( .A(\CACHE[4][145] ), .B(\CACHE[5][145] ), .C(\CACHE[6][145] ), 
        .D(\CACHE[7][145] ), .S0(n422), .S1(n457), .Y(n3387) );
  MXI4X1 U2092 ( .A(\CACHE[0][145] ), .B(\CACHE[1][145] ), .C(\CACHE[2][145] ), 
        .D(\CACHE[3][145] ), .S0(n422), .S1(n457), .Y(n3386) );
  MXI2X1 U2093 ( .A(n3394), .B(n3395), .S0(n470), .Y(N38) );
  MXI4X1 U2094 ( .A(\CACHE[4][149] ), .B(\CACHE[5][149] ), .C(\CACHE[6][149] ), 
        .D(\CACHE[7][149] ), .S0(n431), .S1(n457), .Y(n3395) );
  MXI4X1 U2095 ( .A(\CACHE[0][149] ), .B(\CACHE[1][149] ), .C(\CACHE[2][149] ), 
        .D(\CACHE[3][149] ), .S0(n430), .S1(n457), .Y(n3394) );
  MXI2X1 U2096 ( .A(n3396), .B(n3397), .S0(n470), .Y(N37) );
  MXI4X1 U2097 ( .A(\CACHE[4][150] ), .B(\CACHE[5][150] ), .C(\CACHE[6][150] ), 
        .D(\CACHE[7][150] ), .S0(n428), .S1(n458), .Y(n3397) );
  MXI4X1 U2098 ( .A(\CACHE[0][150] ), .B(\CACHE[1][150] ), .C(\CACHE[2][150] ), 
        .D(\CACHE[3][150] ), .S0(n424), .S1(n458), .Y(n3396) );
  MXI2X1 U2099 ( .A(n3398), .B(n3399), .S0(n470), .Y(N36) );
  MXI4X1 U2100 ( .A(\CACHE[4][151] ), .B(\CACHE[5][151] ), .C(\CACHE[6][151] ), 
        .D(\CACHE[7][151] ), .S0(n433), .S1(n458), .Y(n3399) );
  MXI4X1 U2101 ( .A(\CACHE[0][151] ), .B(\CACHE[1][151] ), .C(\CACHE[2][151] ), 
        .D(\CACHE[3][151] ), .S0(n419), .S1(n458), .Y(n3398) );
  MXI2X1 U2102 ( .A(n3400), .B(n3401), .S0(n470), .Y(N35) );
  MXI4X1 U2103 ( .A(\CACHE[4][152] ), .B(\CACHE[5][152] ), .C(\CACHE[6][152] ), 
        .D(\CACHE[7][152] ), .S0(n418), .S1(n458), .Y(n3401) );
  MXI4X1 U2104 ( .A(\CACHE[0][152] ), .B(\CACHE[1][152] ), .C(\CACHE[2][152] ), 
        .D(\CACHE[3][152] ), .S0(n425), .S1(n458), .Y(n3400) );
  MXI2X1 U2105 ( .A(n3352), .B(n3353), .S0(n468), .Y(N59) );
  MXI4X1 U2106 ( .A(\CACHE[4][128] ), .B(\CACHE[5][128] ), .C(\CACHE[6][128] ), 
        .D(\CACHE[7][128] ), .S0(n419), .S1(n455), .Y(n3353) );
  MXI4X1 U2107 ( .A(\CACHE[0][128] ), .B(\CACHE[1][128] ), .C(\CACHE[2][128] ), 
        .D(\CACHE[3][128] ), .S0(n419), .S1(n455), .Y(n3352) );
  MXI2X1 U2108 ( .A(n3354), .B(n3355), .S0(n468), .Y(N58) );
  MXI4X1 U2109 ( .A(\CACHE[4][129] ), .B(\CACHE[5][129] ), .C(\CACHE[6][129] ), 
        .D(\CACHE[7][129] ), .S0(n419), .S1(n455), .Y(n3355) );
  MXI4X1 U2110 ( .A(\CACHE[0][129] ), .B(\CACHE[1][129] ), .C(\CACHE[2][129] ), 
        .D(\CACHE[3][129] ), .S0(n420), .S1(n455), .Y(n3354) );
  MXI2X1 U2111 ( .A(n3356), .B(n3357), .S0(n468), .Y(N57) );
  MXI4X1 U2112 ( .A(\CACHE[4][130] ), .B(\CACHE[5][130] ), .C(\CACHE[6][130] ), 
        .D(\CACHE[7][130] ), .S0(n420), .S1(n455), .Y(n3357) );
  MXI4X1 U2113 ( .A(\CACHE[0][130] ), .B(\CACHE[1][130] ), .C(\CACHE[2][130] ), 
        .D(\CACHE[3][130] ), .S0(n420), .S1(n455), .Y(n3356) );
  MXI2X1 U2114 ( .A(n3364), .B(n3365), .S0(n469), .Y(N53) );
  MXI4X1 U2115 ( .A(\CACHE[4][134] ), .B(\CACHE[5][134] ), .C(\CACHE[6][134] ), 
        .D(\CACHE[7][134] ), .S0(n420), .S1(n453), .Y(n3365) );
  MXI4X1 U2116 ( .A(\CACHE[0][134] ), .B(\CACHE[1][134] ), .C(\CACHE[2][134] ), 
        .D(\CACHE[3][134] ), .S0(n420), .S1(n444), .Y(n3364) );
  MXI2X1 U2117 ( .A(n3366), .B(n3367), .S0(n469), .Y(N52) );
  MXI4X1 U2118 ( .A(\CACHE[4][135] ), .B(\CACHE[5][135] ), .C(\CACHE[6][135] ), 
        .D(\CACHE[7][135] ), .S0(n420), .S1(n451), .Y(n3367) );
  MXI4X1 U2119 ( .A(\CACHE[0][135] ), .B(\CACHE[1][135] ), .C(\CACHE[2][135] ), 
        .D(\CACHE[3][135] ), .S0(n420), .S1(n455), .Y(n3366) );
  MXI2X1 U2120 ( .A(n3368), .B(n3369), .S0(n469), .Y(N51) );
  MXI4X1 U2121 ( .A(\CACHE[4][136] ), .B(\CACHE[5][136] ), .C(\CACHE[6][136] ), 
        .D(\CACHE[7][136] ), .S0(n421), .S1(n441), .Y(n3369) );
  MXI4X1 U2122 ( .A(\CACHE[0][136] ), .B(\CACHE[1][136] ), .C(\CACHE[2][136] ), 
        .D(\CACHE[3][136] ), .S0(n421), .S1(n457), .Y(n3368) );
  MXI2X1 U2123 ( .A(n3376), .B(n3377), .S0(n469), .Y(N47) );
  MXI4X1 U2124 ( .A(\CACHE[4][140] ), .B(\CACHE[5][140] ), .C(\CACHE[6][140] ), 
        .D(\CACHE[7][140] ), .S0(n421), .S1(n456), .Y(n3377) );
  MXI4X1 U2125 ( .A(\CACHE[0][140] ), .B(\CACHE[1][140] ), .C(\CACHE[2][140] ), 
        .D(\CACHE[3][140] ), .S0(n421), .S1(n456), .Y(n3376) );
  MXI2X1 U2126 ( .A(n3378), .B(n3379), .S0(n469), .Y(N46) );
  MXI4X1 U2127 ( .A(\CACHE[4][141] ), .B(\CACHE[5][141] ), .C(\CACHE[6][141] ), 
        .D(\CACHE[7][141] ), .S0(n421), .S1(n456), .Y(n3379) );
  MXI4X1 U2128 ( .A(\CACHE[0][141] ), .B(\CACHE[1][141] ), .C(\CACHE[2][141] ), 
        .D(\CACHE[3][141] ), .S0(n421), .S1(n456), .Y(n3378) );
  MXI2X1 U2129 ( .A(n3380), .B(n3381), .S0(n469), .Y(N45) );
  MXI4X1 U2130 ( .A(\CACHE[4][142] ), .B(\CACHE[5][142] ), .C(\CACHE[6][142] ), 
        .D(\CACHE[7][142] ), .S0(n421), .S1(n456), .Y(n3381) );
  MXI4X1 U2131 ( .A(\CACHE[0][142] ), .B(\CACHE[1][142] ), .C(\CACHE[2][142] ), 
        .D(\CACHE[3][142] ), .S0(n422), .S1(n456), .Y(n3380) );
  MXI2X1 U2132 ( .A(n3388), .B(n3389), .S0(n470), .Y(N41) );
  MXI4X1 U2133 ( .A(\CACHE[4][146] ), .B(\CACHE[5][146] ), .C(\CACHE[6][146] ), 
        .D(\CACHE[7][146] ), .S0(n422), .S1(n457), .Y(n3389) );
  MXI4X1 U2134 ( .A(\CACHE[0][146] ), .B(\CACHE[1][146] ), .C(\CACHE[2][146] ), 
        .D(\CACHE[3][146] ), .S0(n422), .S1(n457), .Y(n3388) );
  MXI2X1 U2135 ( .A(n3390), .B(n3391), .S0(n470), .Y(N40) );
  MXI4X1 U2136 ( .A(\CACHE[4][147] ), .B(\CACHE[5][147] ), .C(\CACHE[6][147] ), 
        .D(\CACHE[7][147] ), .S0(n422), .S1(n457), .Y(n3391) );
  MXI4X1 U2137 ( .A(\CACHE[0][147] ), .B(\CACHE[1][147] ), .C(\CACHE[2][147] ), 
        .D(\CACHE[3][147] ), .S0(n422), .S1(n457), .Y(n3390) );
  MXI2X1 U2138 ( .A(n3392), .B(n3393), .S0(n470), .Y(N39) );
  MXI4X1 U2139 ( .A(\CACHE[4][148] ), .B(\CACHE[5][148] ), .C(\CACHE[6][148] ), 
        .D(\CACHE[7][148] ), .S0(n422), .S1(n457), .Y(n3393) );
  MXI4X1 U2140 ( .A(\CACHE[0][148] ), .B(\CACHE[1][148] ), .C(\CACHE[2][148] ), 
        .D(\CACHE[3][148] ), .S0(n422), .S1(n457), .Y(n3392) );
  MXI2X1 U2141 ( .A(n3402), .B(n3403), .S0(n470), .Y(N33) );
  MXI4X1 U2142 ( .A(\CACHE[4][154] ), .B(\CACHE[5][154] ), .C(\CACHE[6][154] ), 
        .D(\CACHE[7][154] ), .S0(n429), .S1(n458), .Y(n3403) );
  MXI4X1 U2143 ( .A(\CACHE[0][154] ), .B(\CACHE[1][154] ), .C(\CACHE[2][154] ), 
        .D(\CACHE[3][154] ), .S0(n432), .S1(n458), .Y(n3402) );
  MXI2X1 U2144 ( .A(n3096), .B(n3097), .S0(n462), .Y(N187) );
  MXI4X1 U2145 ( .A(\CACHE[4][0] ), .B(\CACHE[5][0] ), .C(\CACHE[6][0] ), .D(
        \CACHE[7][0] ), .S0(n415), .S1(n438), .Y(n3097) );
  MXI4X1 U2146 ( .A(\CACHE[0][0] ), .B(\CACHE[1][0] ), .C(\CACHE[2][0] ), .D(
        \CACHE[3][0] ), .S0(n428), .S1(n438), .Y(n3096) );
  MXI2X1 U2147 ( .A(n3288), .B(n3289), .S0(n466), .Y(N91) );
  MXI4X1 U2148 ( .A(\CACHE[4][96] ), .B(\CACHE[5][96] ), .C(\CACHE[6][96] ), 
        .D(\CACHE[7][96] ), .S0(n423), .S1(n451), .Y(n3289) );
  MXI4X1 U2149 ( .A(\CACHE[0][96] ), .B(\CACHE[1][96] ), .C(\CACHE[2][96] ), 
        .D(\CACHE[3][96] ), .S0(n417), .S1(n451), .Y(n3288) );
  MXI2X1 U2150 ( .A(n3098), .B(n3099), .S0(n462), .Y(N186) );
  MXI4X1 U2151 ( .A(\CACHE[4][1] ), .B(\CACHE[5][1] ), .C(\CACHE[6][1] ), .D(
        \CACHE[7][1] ), .S0(n423), .S1(n438), .Y(n3099) );
  MXI4X1 U2152 ( .A(\CACHE[0][1] ), .B(\CACHE[1][1] ), .C(\CACHE[2][1] ), .D(
        \CACHE[3][1] ), .S0(n423), .S1(n438), .Y(n3098) );
  MXI2X1 U2153 ( .A(n3290), .B(n3291), .S0(n466), .Y(N90) );
  MXI4X1 U2154 ( .A(\CACHE[4][97] ), .B(\CACHE[5][97] ), .C(\CACHE[6][97] ), 
        .D(\CACHE[7][97] ), .S0(n417), .S1(n451), .Y(n3291) );
  MXI4X1 U2155 ( .A(\CACHE[0][97] ), .B(\CACHE[1][97] ), .C(\CACHE[2][97] ), 
        .D(\CACHE[3][97] ), .S0(n417), .S1(n451), .Y(n3290) );
  MXI2X1 U2156 ( .A(n3100), .B(n3101), .S0(n462), .Y(N185) );
  MXI4X1 U2157 ( .A(\CACHE[4][2] ), .B(\CACHE[5][2] ), .C(\CACHE[6][2] ), .D(
        \CACHE[7][2] ), .S0(n423), .S1(n438), .Y(n3101) );
  MXI4X1 U2158 ( .A(\CACHE[0][2] ), .B(\CACHE[1][2] ), .C(\CACHE[2][2] ), .D(
        \CACHE[3][2] ), .S0(n423), .S1(n438), .Y(n3100) );
  MXI2X1 U2159 ( .A(n3292), .B(n3293), .S0(n466), .Y(N89) );
  MXI4X1 U2160 ( .A(\CACHE[4][98] ), .B(\CACHE[5][98] ), .C(\CACHE[6][98] ), 
        .D(\CACHE[7][98] ), .S0(n417), .S1(n451), .Y(n3293) );
  MXI4X1 U2161 ( .A(\CACHE[0][98] ), .B(\CACHE[1][98] ), .C(\CACHE[2][98] ), 
        .D(\CACHE[3][98] ), .S0(n417), .S1(n451), .Y(n3292) );
  MXI2X1 U2162 ( .A(n3102), .B(n3103), .S0(n462), .Y(N184) );
  MXI4X1 U2163 ( .A(\CACHE[4][3] ), .B(\CACHE[5][3] ), .C(\CACHE[6][3] ), .D(
        \CACHE[7][3] ), .S0(n423), .S1(n438), .Y(n3103) );
  MXI4X1 U2164 ( .A(\CACHE[0][3] ), .B(\CACHE[1][3] ), .C(\CACHE[2][3] ), .D(
        \CACHE[3][3] ), .S0(n423), .S1(n438), .Y(n3102) );
  MXI2X1 U2165 ( .A(n3294), .B(n3295), .S0(n466), .Y(N88) );
  MXI4X1 U2166 ( .A(\CACHE[4][99] ), .B(\CACHE[5][99] ), .C(\CACHE[6][99] ), 
        .D(\CACHE[7][99] ), .S0(n417), .S1(n451), .Y(n3295) );
  MXI4X1 U2167 ( .A(\CACHE[0][99] ), .B(\CACHE[1][99] ), .C(\CACHE[2][99] ), 
        .D(\CACHE[3][99] ), .S0(n417), .S1(n451), .Y(n3294) );
  MXI2X1 U2168 ( .A(n3104), .B(n3105), .S0(n462), .Y(N183) );
  MXI4X1 U2169 ( .A(\CACHE[4][4] ), .B(\CACHE[5][4] ), .C(\CACHE[6][4] ), .D(
        \CACHE[7][4] ), .S0(n423), .S1(n438), .Y(n3105) );
  MXI4X1 U2170 ( .A(\CACHE[0][4] ), .B(\CACHE[1][4] ), .C(\CACHE[2][4] ), .D(
        \CACHE[3][4] ), .S0(n423), .S1(n438), .Y(n3104) );
  MXI2X1 U2171 ( .A(n3296), .B(n3297), .S0(n466), .Y(N87) );
  MXI4X1 U2172 ( .A(\CACHE[4][100] ), .B(\CACHE[5][100] ), .C(\CACHE[6][100] ), 
        .D(\CACHE[7][100] ), .S0(n417), .S1(n451), .Y(n3297) );
  MXI4X1 U2173 ( .A(\CACHE[0][100] ), .B(\CACHE[1][100] ), .C(\CACHE[2][100] ), 
        .D(\CACHE[3][100] ), .S0(n417), .S1(n451), .Y(n3296) );
  MXI2X1 U2174 ( .A(n3106), .B(n3107), .S0(n462), .Y(N182) );
  MXI4X1 U2175 ( .A(\CACHE[4][5] ), .B(\CACHE[5][5] ), .C(\CACHE[6][5] ), .D(
        \CACHE[7][5] ), .S0(n423), .S1(n438), .Y(n3107) );
  MXI4X1 U2176 ( .A(\CACHE[0][5] ), .B(\CACHE[1][5] ), .C(\CACHE[2][5] ), .D(
        \CACHE[3][5] ), .S0(n423), .S1(n438), .Y(n3106) );
  MXI2X1 U2177 ( .A(n3298), .B(n3299), .S0(n466), .Y(N86) );
  MXI4X1 U2178 ( .A(\CACHE[4][101] ), .B(\CACHE[5][101] ), .C(\CACHE[6][101] ), 
        .D(\CACHE[7][101] ), .S0(n417), .S1(n451), .Y(n3299) );
  MXI4X1 U2179 ( .A(\CACHE[0][101] ), .B(\CACHE[1][101] ), .C(\CACHE[2][101] ), 
        .D(\CACHE[3][101] ), .S0(n417), .S1(n451), .Y(n3298) );
  MXI2X1 U2180 ( .A(n3108), .B(n3109), .S0(n462), .Y(N181) );
  MXI4X1 U2181 ( .A(\CACHE[4][6] ), .B(\CACHE[5][6] ), .C(\CACHE[6][6] ), .D(
        \CACHE[7][6] ), .S0(n423), .S1(n439), .Y(n3109) );
  MXI4X1 U2182 ( .A(\CACHE[0][6] ), .B(\CACHE[1][6] ), .C(\CACHE[2][6] ), .D(
        \CACHE[3][6] ), .S0(n423), .S1(n439), .Y(n3108) );
  MXI2X1 U2183 ( .A(n3300), .B(n3301), .S0(n466), .Y(N85) );
  MXI4X1 U2184 ( .A(\CACHE[4][102] ), .B(\CACHE[5][102] ), .C(\CACHE[6][102] ), 
        .D(\CACHE[7][102] ), .S0(n417), .S1(n452), .Y(n3301) );
  MXI4X1 U2185 ( .A(\CACHE[0][102] ), .B(\CACHE[1][102] ), .C(\CACHE[2][102] ), 
        .D(\CACHE[3][102] ), .S0(n417), .S1(n452), .Y(n3300) );
  MXI2X1 U2186 ( .A(n3110), .B(n3111), .S0(n462), .Y(N180) );
  MXI4X1 U2187 ( .A(\CACHE[4][7] ), .B(\CACHE[5][7] ), .C(\CACHE[6][7] ), .D(
        \CACHE[7][7] ), .S0(n423), .S1(n439), .Y(n3111) );
  MXI4X1 U2188 ( .A(\CACHE[0][7] ), .B(\CACHE[1][7] ), .C(\CACHE[2][7] ), .D(
        \CACHE[3][7] ), .S0(n424), .S1(n439), .Y(n3110) );
  MXI2X1 U2189 ( .A(n3302), .B(n3303), .S0(n466), .Y(N84) );
  MXI4X1 U2190 ( .A(\CACHE[4][103] ), .B(\CACHE[5][103] ), .C(\CACHE[6][103] ), 
        .D(\CACHE[7][103] ), .S0(n417), .S1(n452), .Y(n3303) );
  MXI4X1 U2191 ( .A(\CACHE[0][103] ), .B(\CACHE[1][103] ), .C(\CACHE[2][103] ), 
        .D(\CACHE[3][103] ), .S0(n418), .S1(n452), .Y(n3302) );
  MXI2X1 U2192 ( .A(n3112), .B(n3113), .S0(n462), .Y(N179) );
  MXI4X1 U2193 ( .A(\CACHE[4][8] ), .B(\CACHE[5][8] ), .C(\CACHE[6][8] ), .D(
        \CACHE[7][8] ), .S0(n424), .S1(n439), .Y(n3113) );
  MXI4X1 U2194 ( .A(\CACHE[0][8] ), .B(\CACHE[1][8] ), .C(\CACHE[2][8] ), .D(
        \CACHE[3][8] ), .S0(n424), .S1(n439), .Y(n3112) );
  MXI2X1 U2195 ( .A(n3304), .B(n3305), .S0(n466), .Y(N83) );
  MXI4X1 U2196 ( .A(\CACHE[4][104] ), .B(\CACHE[5][104] ), .C(\CACHE[6][104] ), 
        .D(\CACHE[7][104] ), .S0(n418), .S1(n452), .Y(n3305) );
  MXI4X1 U2197 ( .A(\CACHE[0][104] ), .B(\CACHE[1][104] ), .C(\CACHE[2][104] ), 
        .D(\CACHE[3][104] ), .S0(n418), .S1(n452), .Y(n3304) );
  MXI2X1 U2198 ( .A(n3114), .B(n3115), .S0(n462), .Y(N178) );
  MXI4X1 U2199 ( .A(\CACHE[4][9] ), .B(\CACHE[5][9] ), .C(\CACHE[6][9] ), .D(
        \CACHE[7][9] ), .S0(n424), .S1(n439), .Y(n3115) );
  MXI4X1 U2200 ( .A(\CACHE[0][9] ), .B(\CACHE[1][9] ), .C(\CACHE[2][9] ), .D(
        \CACHE[3][9] ), .S0(n424), .S1(n439), .Y(n3114) );
  MXI2X1 U2201 ( .A(n3306), .B(n3307), .S0(n466), .Y(N82) );
  MXI4X1 U2202 ( .A(\CACHE[4][105] ), .B(\CACHE[5][105] ), .C(\CACHE[6][105] ), 
        .D(\CACHE[7][105] ), .S0(n418), .S1(n452), .Y(n3307) );
  MXI4X1 U2203 ( .A(\CACHE[0][105] ), .B(\CACHE[1][105] ), .C(\CACHE[2][105] ), 
        .D(\CACHE[3][105] ), .S0(n418), .S1(n452), .Y(n3306) );
  MXI2X1 U2204 ( .A(n3116), .B(n3117), .S0(n462), .Y(N177) );
  MXI4X1 U2205 ( .A(\CACHE[4][10] ), .B(\CACHE[5][10] ), .C(\CACHE[6][10] ), 
        .D(\CACHE[7][10] ), .S0(n424), .S1(n439), .Y(n3117) );
  MXI4X1 U2206 ( .A(\CACHE[0][10] ), .B(\CACHE[1][10] ), .C(\CACHE[2][10] ), 
        .D(\CACHE[3][10] ), .S0(n424), .S1(n439), .Y(n3116) );
  MXI2X1 U2207 ( .A(n3308), .B(n3309), .S0(n466), .Y(N81) );
  MXI4X1 U2208 ( .A(\CACHE[4][106] ), .B(\CACHE[5][106] ), .C(\CACHE[6][106] ), 
        .D(\CACHE[7][106] ), .S0(n418), .S1(n452), .Y(n3309) );
  MXI4X1 U2209 ( .A(\CACHE[0][106] ), .B(\CACHE[1][106] ), .C(\CACHE[2][106] ), 
        .D(\CACHE[3][106] ), .S0(n418), .S1(n452), .Y(n3308) );
  MXI2X1 U2210 ( .A(n3118), .B(n3119), .S0(n462), .Y(N176) );
  MXI4X1 U2211 ( .A(\CACHE[4][11] ), .B(\CACHE[5][11] ), .C(\CACHE[6][11] ), 
        .D(\CACHE[7][11] ), .S0(n424), .S1(n439), .Y(n3119) );
  MXI4X1 U2212 ( .A(\CACHE[0][11] ), .B(\CACHE[1][11] ), .C(\CACHE[2][11] ), 
        .D(\CACHE[3][11] ), .S0(n424), .S1(n439), .Y(n3118) );
  MXI2X1 U2213 ( .A(n3310), .B(n3311), .S0(n466), .Y(N80) );
  MXI4X1 U2214 ( .A(\CACHE[4][107] ), .B(\CACHE[5][107] ), .C(\CACHE[6][107] ), 
        .D(\CACHE[7][107] ), .S0(n418), .S1(n452), .Y(n3311) );
  MXI4X1 U2215 ( .A(\CACHE[0][107] ), .B(\CACHE[1][107] ), .C(\CACHE[2][107] ), 
        .D(\CACHE[3][107] ), .S0(n418), .S1(n452), .Y(n3310) );
  MXI2X1 U2216 ( .A(n3120), .B(n3121), .S0(n463), .Y(N175) );
  MXI4X1 U2217 ( .A(\CACHE[4][12] ), .B(\CACHE[5][12] ), .C(\CACHE[6][12] ), 
        .D(\CACHE[7][12] ), .S0(n424), .S1(n440), .Y(n3121) );
  MXI4X1 U2218 ( .A(\CACHE[0][12] ), .B(\CACHE[1][12] ), .C(\CACHE[2][12] ), 
        .D(\CACHE[3][12] ), .S0(n424), .S1(n440), .Y(n3120) );
  MXI2X1 U2219 ( .A(n3312), .B(n3313), .S0(n467), .Y(N79) );
  MXI4X1 U2220 ( .A(\CACHE[4][108] ), .B(\CACHE[5][108] ), .C(\CACHE[6][108] ), 
        .D(\CACHE[7][108] ), .S0(n418), .S1(n453), .Y(n3313) );
  MXI4X1 U2221 ( .A(\CACHE[0][108] ), .B(\CACHE[1][108] ), .C(\CACHE[2][108] ), 
        .D(\CACHE[3][108] ), .S0(n418), .S1(n453), .Y(n3312) );
  MXI2X1 U2222 ( .A(n3122), .B(n3123), .S0(n463), .Y(N174) );
  MXI4X1 U2223 ( .A(\CACHE[4][13] ), .B(\CACHE[5][13] ), .C(\CACHE[6][13] ), 
        .D(\CACHE[7][13] ), .S0(n424), .S1(n440), .Y(n3123) );
  MXI4X1 U2224 ( .A(\CACHE[0][13] ), .B(\CACHE[1][13] ), .C(\CACHE[2][13] ), 
        .D(\CACHE[3][13] ), .S0(n424), .S1(n440), .Y(n3122) );
  MXI2X1 U2225 ( .A(n3314), .B(n3315), .S0(n467), .Y(N78) );
  MXI4X1 U2226 ( .A(\CACHE[4][109] ), .B(\CACHE[5][109] ), .C(\CACHE[6][109] ), 
        .D(\CACHE[7][109] ), .S0(n418), .S1(n453), .Y(n3315) );
  MXI4X1 U2227 ( .A(\CACHE[0][109] ), .B(\CACHE[1][109] ), .C(\CACHE[2][109] ), 
        .D(\CACHE[3][109] ), .S0(n418), .S1(n453), .Y(n3314) );
  MXI2X1 U2228 ( .A(n3124), .B(n3125), .S0(n463), .Y(N173) );
  MXI4X1 U2229 ( .A(\CACHE[4][14] ), .B(\CACHE[5][14] ), .C(\CACHE[6][14] ), 
        .D(\CACHE[7][14] ), .S0(n425), .S1(n440), .Y(n3125) );
  MXI4X1 U2230 ( .A(\CACHE[0][14] ), .B(\CACHE[1][14] ), .C(\CACHE[2][14] ), 
        .D(\CACHE[3][14] ), .S0(n425), .S1(n440), .Y(n3124) );
  MXI2X1 U2231 ( .A(n3316), .B(n3317), .S0(n467), .Y(N77) );
  MXI4X1 U2232 ( .A(\CACHE[4][110] ), .B(\CACHE[5][110] ), .C(\CACHE[6][110] ), 
        .D(\CACHE[7][110] ), .S0(n419), .S1(n453), .Y(n3317) );
  MXI4X1 U2233 ( .A(\CACHE[0][110] ), .B(\CACHE[1][110] ), .C(\CACHE[2][110] ), 
        .D(\CACHE[3][110] ), .S0(n428), .S1(n453), .Y(n3316) );
  MXI2X1 U2234 ( .A(n3126), .B(n3127), .S0(n463), .Y(N172) );
  MXI4X1 U2235 ( .A(\CACHE[4][15] ), .B(\CACHE[5][15] ), .C(\CACHE[6][15] ), 
        .D(\CACHE[7][15] ), .S0(n425), .S1(n440), .Y(n3127) );
  MXI4X1 U2236 ( .A(\CACHE[0][15] ), .B(\CACHE[1][15] ), .C(\CACHE[2][15] ), 
        .D(\CACHE[3][15] ), .S0(n425), .S1(n440), .Y(n3126) );
  MXI2X1 U2237 ( .A(n3318), .B(n3319), .S0(n467), .Y(N76) );
  MXI4X1 U2238 ( .A(\CACHE[4][111] ), .B(\CACHE[5][111] ), .C(\CACHE[6][111] ), 
        .D(\CACHE[7][111] ), .S0(n432), .S1(n453), .Y(n3319) );
  MXI4X1 U2239 ( .A(\CACHE[0][111] ), .B(\CACHE[1][111] ), .C(\CACHE[2][111] ), 
        .D(\CACHE[3][111] ), .S0(n418), .S1(n453), .Y(n3318) );
  MXI2X1 U2240 ( .A(n3128), .B(n3129), .S0(n463), .Y(N171) );
  MXI4X1 U2241 ( .A(\CACHE[4][16] ), .B(\CACHE[5][16] ), .C(\CACHE[6][16] ), 
        .D(\CACHE[7][16] ), .S0(n425), .S1(n440), .Y(n3129) );
  MXI4X1 U2242 ( .A(\CACHE[0][16] ), .B(\CACHE[1][16] ), .C(\CACHE[2][16] ), 
        .D(\CACHE[3][16] ), .S0(n425), .S1(n440), .Y(n3128) );
  MXI2X1 U2243 ( .A(n3320), .B(n3321), .S0(n467), .Y(N75) );
  MXI4X1 U2244 ( .A(\CACHE[4][112] ), .B(\CACHE[5][112] ), .C(\CACHE[6][112] ), 
        .D(\CACHE[7][112] ), .S0(n415), .S1(n453), .Y(n3321) );
  MXI4X1 U2245 ( .A(\CACHE[0][112] ), .B(\CACHE[1][112] ), .C(\CACHE[2][112] ), 
        .D(\CACHE[3][112] ), .S0(n429), .S1(n453), .Y(n3320) );
  MXI2X1 U2246 ( .A(n3130), .B(n3131), .S0(n463), .Y(N170) );
  MXI4X1 U2247 ( .A(\CACHE[4][17] ), .B(\CACHE[5][17] ), .C(\CACHE[6][17] ), 
        .D(\CACHE[7][17] ), .S0(n425), .S1(n440), .Y(n3131) );
  MXI4X1 U2248 ( .A(\CACHE[0][17] ), .B(\CACHE[1][17] ), .C(\CACHE[2][17] ), 
        .D(\CACHE[3][17] ), .S0(n425), .S1(n440), .Y(n3130) );
  MXI2X1 U2249 ( .A(n3322), .B(n3323), .S0(n467), .Y(N74) );
  MXI4X1 U2250 ( .A(\CACHE[4][113] ), .B(\CACHE[5][113] ), .C(\CACHE[6][113] ), 
        .D(\CACHE[7][113] ), .S0(n427), .S1(n453), .Y(n3323) );
  MXI4X1 U2251 ( .A(\CACHE[0][113] ), .B(\CACHE[1][113] ), .C(\CACHE[2][113] ), 
        .D(\CACHE[3][113] ), .S0(n416), .S1(n453), .Y(n3322) );
  MXI2X1 U2252 ( .A(n3132), .B(n3133), .S0(n463), .Y(N169) );
  MXI4X1 U2253 ( .A(\CACHE[4][18] ), .B(\CACHE[5][18] ), .C(\CACHE[6][18] ), 
        .D(\CACHE[7][18] ), .S0(n425), .S1(n441), .Y(n3133) );
  MXI4X1 U2254 ( .A(\CACHE[0][18] ), .B(\CACHE[1][18] ), .C(\CACHE[2][18] ), 
        .D(\CACHE[3][18] ), .S0(n425), .S1(n441), .Y(n3132) );
  MXI2X1 U2255 ( .A(n3324), .B(n3325), .S0(n467), .Y(N73) );
  MXI4X1 U2256 ( .A(\CACHE[4][114] ), .B(\CACHE[5][114] ), .C(\CACHE[6][114] ), 
        .D(\CACHE[7][114] ), .S0(n420), .S1(n454), .Y(n3325) );
  MXI4X1 U2257 ( .A(\CACHE[0][114] ), .B(\CACHE[1][114] ), .C(\CACHE[2][114] ), 
        .D(\CACHE[3][114] ), .S0(n430), .S1(n454), .Y(n3324) );
  MXI2X1 U2258 ( .A(n3134), .B(n3135), .S0(n463), .Y(N168) );
  MXI4X1 U2259 ( .A(\CACHE[4][19] ), .B(\CACHE[5][19] ), .C(\CACHE[6][19] ), 
        .D(\CACHE[7][19] ), .S0(n425), .S1(n441), .Y(n3135) );
  MXI4X1 U2260 ( .A(\CACHE[0][19] ), .B(\CACHE[1][19] ), .C(\CACHE[2][19] ), 
        .D(\CACHE[3][19] ), .S0(n425), .S1(n441), .Y(n3134) );
  MXI2X1 U2261 ( .A(n3326), .B(n3327), .S0(n467), .Y(N72) );
  MXI4X1 U2262 ( .A(\CACHE[4][115] ), .B(\CACHE[5][115] ), .C(\CACHE[6][115] ), 
        .D(\CACHE[7][115] ), .S0(n422), .S1(n454), .Y(n3327) );
  MXI4X1 U2263 ( .A(\CACHE[0][115] ), .B(\CACHE[1][115] ), .C(\CACHE[2][115] ), 
        .D(\CACHE[3][115] ), .S0(n417), .S1(n454), .Y(n3326) );
  MXI2X1 U2264 ( .A(n3136), .B(n3137), .S0(n463), .Y(N167) );
  MXI4X1 U2265 ( .A(\CACHE[4][20] ), .B(\CACHE[5][20] ), .C(\CACHE[6][20] ), 
        .D(\CACHE[7][20] ), .S0(n425), .S1(n441), .Y(n3137) );
  MXI4X1 U2266 ( .A(\CACHE[0][20] ), .B(\CACHE[1][20] ), .C(\CACHE[2][20] ), 
        .D(\CACHE[3][20] ), .S0(n426), .S1(n441), .Y(n3136) );
  MXI2X1 U2267 ( .A(n3328), .B(n3329), .S0(n467), .Y(N71) );
  MXI4X1 U2268 ( .A(\CACHE[4][116] ), .B(\CACHE[5][116] ), .C(\CACHE[6][116] ), 
        .D(\CACHE[7][116] ), .S0(n424), .S1(n454), .Y(n3329) );
  MXI4X1 U2269 ( .A(\CACHE[0][116] ), .B(\CACHE[1][116] ), .C(\CACHE[2][116] ), 
        .D(\CACHE[3][116] ), .S0(n431), .S1(n454), .Y(n3328) );
  MXI2X1 U2270 ( .A(n3138), .B(n3139), .S0(n463), .Y(N166) );
  MXI4X1 U2271 ( .A(\CACHE[4][21] ), .B(\CACHE[5][21] ), .C(\CACHE[6][21] ), 
        .D(\CACHE[7][21] ), .S0(n426), .S1(n441), .Y(n3139) );
  MXI4X1 U2272 ( .A(\CACHE[0][21] ), .B(\CACHE[1][21] ), .C(\CACHE[2][21] ), 
        .D(\CACHE[3][21] ), .S0(n426), .S1(n441), .Y(n3138) );
  MXI2X1 U2273 ( .A(n3330), .B(n3331), .S0(n467), .Y(N70) );
  MXI4X1 U2274 ( .A(\CACHE[4][117] ), .B(\CACHE[5][117] ), .C(\CACHE[6][117] ), 
        .D(\CACHE[7][117] ), .S0(n428), .S1(n454), .Y(n3331) );
  MXI4X1 U2275 ( .A(\CACHE[0][117] ), .B(\CACHE[1][117] ), .C(\CACHE[2][117] ), 
        .D(\CACHE[3][117] ), .S0(n415), .S1(n454), .Y(n3330) );
  MXI2X1 U2276 ( .A(n3140), .B(n3141), .S0(n463), .Y(N165) );
  MXI4X1 U2277 ( .A(\CACHE[4][22] ), .B(\CACHE[5][22] ), .C(\CACHE[6][22] ), 
        .D(\CACHE[7][22] ), .S0(n426), .S1(n441), .Y(n3141) );
  MXI4X1 U2278 ( .A(\CACHE[0][22] ), .B(\CACHE[1][22] ), .C(\CACHE[2][22] ), 
        .D(\CACHE[3][22] ), .S0(n426), .S1(n441), .Y(n3140) );
  MXI2X1 U2279 ( .A(n3332), .B(n3333), .S0(n467), .Y(N69) );
  MXI4X1 U2280 ( .A(\CACHE[4][118] ), .B(\CACHE[5][118] ), .C(\CACHE[6][118] ), 
        .D(\CACHE[7][118] ), .S0(n433), .S1(n454), .Y(n3333) );
  MXI4X1 U2281 ( .A(\CACHE[0][118] ), .B(\CACHE[1][118] ), .C(\CACHE[2][118] ), 
        .D(\CACHE[3][118] ), .S0(n419), .S1(n454), .Y(n3332) );
  MXI2X1 U2282 ( .A(n3142), .B(n3143), .S0(n463), .Y(N164) );
  MXI4X1 U2283 ( .A(\CACHE[4][23] ), .B(\CACHE[5][23] ), .C(\CACHE[6][23] ), 
        .D(\CACHE[7][23] ), .S0(n426), .S1(n441), .Y(n3143) );
  MXI4X1 U2284 ( .A(\CACHE[0][23] ), .B(\CACHE[1][23] ), .C(\CACHE[2][23] ), 
        .D(\CACHE[3][23] ), .S0(n426), .S1(n441), .Y(n3142) );
  MXI2X1 U2285 ( .A(n3334), .B(n3335), .S0(n467), .Y(N68) );
  MXI4X1 U2286 ( .A(\CACHE[4][119] ), .B(\CACHE[5][119] ), .C(\CACHE[6][119] ), 
        .D(\CACHE[7][119] ), .S0(n418), .S1(n454), .Y(n3335) );
  MXI4X1 U2287 ( .A(\CACHE[0][119] ), .B(\CACHE[1][119] ), .C(\CACHE[2][119] ), 
        .D(\CACHE[3][119] ), .S0(n425), .S1(n454), .Y(n3334) );
  MXI2X1 U2288 ( .A(n3144), .B(n3145), .S0(n464), .Y(N163) );
  MXI4X1 U2289 ( .A(\CACHE[4][24] ), .B(\CACHE[5][24] ), .C(\CACHE[6][24] ), 
        .D(\CACHE[7][24] ), .S0(n426), .S1(n442), .Y(n3145) );
  MXI4X1 U2290 ( .A(\CACHE[0][24] ), .B(\CACHE[1][24] ), .C(\CACHE[2][24] ), 
        .D(\CACHE[3][24] ), .S0(n426), .S1(n442), .Y(n3144) );
  MXI2X1 U2291 ( .A(n3336), .B(n3337), .S0(n468), .Y(N67) );
  MXI4X1 U2292 ( .A(\CACHE[4][120] ), .B(\CACHE[5][120] ), .C(\CACHE[6][120] ), 
        .D(\CACHE[7][120] ), .S0(n429), .S1(n449), .Y(n3337) );
  MXI4X1 U2293 ( .A(\CACHE[0][120] ), .B(\CACHE[1][120] ), .C(\CACHE[2][120] ), 
        .D(\CACHE[3][120] ), .S0(n432), .S1(n454), .Y(n3336) );
  MXI2X1 U2294 ( .A(n3146), .B(n3147), .S0(n464), .Y(N162) );
  MXI4X1 U2295 ( .A(\CACHE[4][25] ), .B(\CACHE[5][25] ), .C(\CACHE[6][25] ), 
        .D(\CACHE[7][25] ), .S0(n426), .S1(n442), .Y(n3147) );
  MXI4X1 U2296 ( .A(\CACHE[0][25] ), .B(\CACHE[1][25] ), .C(\CACHE[2][25] ), 
        .D(\CACHE[3][25] ), .S0(n426), .S1(n442), .Y(n3146) );
  MXI2X1 U2297 ( .A(n3338), .B(n3339), .S0(n468), .Y(N66) );
  MXI4X1 U2298 ( .A(\CACHE[4][121] ), .B(\CACHE[5][121] ), .C(\CACHE[6][121] ), 
        .D(\CACHE[7][121] ), .S0(n416), .S1(n446), .Y(n3339) );
  MXI4X1 U2299 ( .A(\CACHE[0][121] ), .B(\CACHE[1][121] ), .C(\CACHE[2][121] ), 
        .D(\CACHE[3][121] ), .S0(n415), .S1(n445), .Y(n3338) );
  MXI2X1 U2300 ( .A(n3148), .B(n3149), .S0(n464), .Y(N161) );
  MXI4X1 U2301 ( .A(\CACHE[4][26] ), .B(\CACHE[5][26] ), .C(\CACHE[6][26] ), 
        .D(\CACHE[7][26] ), .S0(n426), .S1(n442), .Y(n3149) );
  MXI4X1 U2302 ( .A(\CACHE[0][26] ), .B(\CACHE[1][26] ), .C(\CACHE[2][26] ), 
        .D(\CACHE[3][26] ), .S0(n426), .S1(n442), .Y(n3148) );
  MXI2X1 U2303 ( .A(n3340), .B(n3341), .S0(n468), .Y(N65) );
  MXI4X1 U2304 ( .A(\CACHE[4][122] ), .B(\CACHE[5][122] ), .C(\CACHE[6][122] ), 
        .D(\CACHE[7][122] ), .S0(n420), .S1(n458), .Y(n3341) );
  MXI4X1 U2305 ( .A(\CACHE[0][122] ), .B(\CACHE[1][122] ), .C(\CACHE[2][122] ), 
        .D(\CACHE[3][122] ), .S0(n427), .S1(n447), .Y(n3340) );
  MXI2X1 U2306 ( .A(n3150), .B(n3151), .S0(n464), .Y(N160) );
  MXI4X1 U2307 ( .A(\CACHE[4][27] ), .B(\CACHE[5][27] ), .C(\CACHE[6][27] ), 
        .D(\CACHE[7][27] ), .S0(n427), .S1(n442), .Y(n3151) );
  MXI4X1 U2308 ( .A(\CACHE[0][27] ), .B(\CACHE[1][27] ), .C(\CACHE[2][27] ), 
        .D(\CACHE[3][27] ), .S0(n427), .S1(n442), .Y(n3150) );
  MXI2X1 U2309 ( .A(n3342), .B(n3343), .S0(n468), .Y(N64) );
  MXI4X1 U2310 ( .A(\CACHE[4][123] ), .B(\CACHE[5][123] ), .C(\CACHE[6][123] ), 
        .D(\CACHE[7][123] ), .S0(n419), .S1(n450), .Y(n3343) );
  MXI4X1 U2311 ( .A(\CACHE[0][123] ), .B(\CACHE[1][123] ), .C(\CACHE[2][123] ), 
        .D(\CACHE[3][123] ), .S0(n419), .S1(n452), .Y(n3342) );
  MXI2X1 U2312 ( .A(n3152), .B(n3153), .S0(n464), .Y(N159) );
  MXI4X1 U2313 ( .A(\CACHE[4][28] ), .B(\CACHE[5][28] ), .C(\CACHE[6][28] ), 
        .D(\CACHE[7][28] ), .S0(n427), .S1(n442), .Y(n3153) );
  MXI4X1 U2314 ( .A(\CACHE[0][28] ), .B(\CACHE[1][28] ), .C(\CACHE[2][28] ), 
        .D(\CACHE[3][28] ), .S0(n427), .S1(n442), .Y(n3152) );
  MXI2X1 U2315 ( .A(n3344), .B(n3345), .S0(n468), .Y(N63) );
  MXI4X1 U2316 ( .A(\CACHE[4][124] ), .B(\CACHE[5][124] ), .C(\CACHE[6][124] ), 
        .D(\CACHE[7][124] ), .S0(n419), .S1(n438), .Y(n3345) );
  MXI4X1 U2317 ( .A(\CACHE[0][124] ), .B(\CACHE[1][124] ), .C(\CACHE[2][124] ), 
        .D(\CACHE[3][124] ), .S0(n419), .S1(n443), .Y(n3344) );
  MXI2X1 U2318 ( .A(n3154), .B(n3155), .S0(n464), .Y(N158) );
  MXI4X1 U2319 ( .A(\CACHE[4][29] ), .B(\CACHE[5][29] ), .C(\CACHE[6][29] ), 
        .D(\CACHE[7][29] ), .S0(n427), .S1(n442), .Y(n3155) );
  MXI4X1 U2320 ( .A(\CACHE[0][29] ), .B(\CACHE[1][29] ), .C(\CACHE[2][29] ), 
        .D(\CACHE[3][29] ), .S0(n427), .S1(n442), .Y(n3154) );
  MXI2X1 U2321 ( .A(n3346), .B(n3347), .S0(n468), .Y(N62) );
  MXI4X1 U2322 ( .A(\CACHE[4][125] ), .B(\CACHE[5][125] ), .C(\CACHE[6][125] ), 
        .D(\CACHE[7][125] ), .S0(n419), .S1(n448), .Y(n3347) );
  MXI4X1 U2323 ( .A(\CACHE[0][125] ), .B(\CACHE[1][125] ), .C(\CACHE[2][125] ), 
        .D(\CACHE[3][125] ), .S0(n419), .S1(n440), .Y(n3346) );
  MXI2X1 U2324 ( .A(n3156), .B(n3157), .S0(n464), .Y(N157) );
  MXI4X1 U2325 ( .A(\CACHE[4][30] ), .B(\CACHE[5][30] ), .C(\CACHE[6][30] ), 
        .D(\CACHE[7][30] ), .S0(n427), .S1(n438), .Y(n3157) );
  MXI4X1 U2326 ( .A(\CACHE[0][30] ), .B(\CACHE[1][30] ), .C(\CACHE[2][30] ), 
        .D(\CACHE[3][30] ), .S0(n427), .S1(n443), .Y(n3156) );
  MXI2X1 U2327 ( .A(n3348), .B(n3349), .S0(n468), .Y(N61) );
  MXI4X1 U2328 ( .A(\CACHE[4][126] ), .B(\CACHE[5][126] ), .C(\CACHE[6][126] ), 
        .D(\CACHE[7][126] ), .S0(n419), .S1(n455), .Y(n3349) );
  MXI4X1 U2329 ( .A(\CACHE[0][126] ), .B(\CACHE[1][126] ), .C(\CACHE[2][126] ), 
        .D(\CACHE[3][126] ), .S0(n419), .S1(n455), .Y(n3348) );
  MXI2X1 U2330 ( .A(n3158), .B(n3159), .S0(n464), .Y(N156) );
  MXI4X1 U2331 ( .A(\CACHE[4][31] ), .B(\CACHE[5][31] ), .C(\CACHE[6][31] ), 
        .D(\CACHE[7][31] ), .S0(n427), .S1(n454), .Y(n3159) );
  MXI4X1 U2332 ( .A(\CACHE[0][31] ), .B(\CACHE[1][31] ), .C(\CACHE[2][31] ), 
        .D(\CACHE[3][31] ), .S0(n427), .S1(n440), .Y(n3158) );
  MXI2X1 U2333 ( .A(n3350), .B(n3351), .S0(n468), .Y(N60) );
  MXI4X1 U2334 ( .A(\CACHE[4][127] ), .B(\CACHE[5][127] ), .C(\CACHE[6][127] ), 
        .D(\CACHE[7][127] ), .S0(n419), .S1(n455), .Y(n3351) );
  MXI4X1 U2335 ( .A(\CACHE[0][127] ), .B(\CACHE[1][127] ), .C(\CACHE[2][127] ), 
        .D(\CACHE[3][127] ), .S0(n419), .S1(n455), .Y(n3350) );
  MXI2X1 U2336 ( .A(n3160), .B(n3161), .S0(n464), .Y(N155) );
  MXI4X1 U2337 ( .A(\CACHE[4][32] ), .B(\CACHE[5][32] ), .C(\CACHE[6][32] ), 
        .D(\CACHE[7][32] ), .S0(n427), .S1(n445), .Y(n3161) );
  MXI4X1 U2338 ( .A(\CACHE[0][32] ), .B(\CACHE[1][32] ), .C(\CACHE[2][32] ), 
        .D(\CACHE[3][32] ), .S0(n427), .S1(n449), .Y(n3160) );
  MXI2X1 U2339 ( .A(n3162), .B(n3163), .S0(n464), .Y(N154) );
  MXI4X1 U2340 ( .A(\CACHE[4][33] ), .B(\CACHE[5][33] ), .C(\CACHE[6][33] ), 
        .D(\CACHE[7][33] ), .S0(n427), .S1(n447), .Y(n3163) );
  MXI4X1 U2341 ( .A(\CACHE[0][33] ), .B(\CACHE[1][33] ), .C(\CACHE[2][33] ), 
        .D(\CACHE[3][33] ), .S0(n428), .S1(n446), .Y(n3162) );
  MXI2X1 U2342 ( .A(n3164), .B(n3165), .S0(n464), .Y(N153) );
  MXI4X1 U2343 ( .A(\CACHE[4][34] ), .B(\CACHE[5][34] ), .C(\CACHE[6][34] ), 
        .D(\CACHE[7][34] ), .S0(n428), .S1(n439), .Y(n3165) );
  MXI4X1 U2344 ( .A(\CACHE[0][34] ), .B(\CACHE[1][34] ), .C(\CACHE[2][34] ), 
        .D(\CACHE[3][34] ), .S0(n428), .S1(n456), .Y(n3164) );
  MXI2X1 U2345 ( .A(n3166), .B(n3167), .S0(n464), .Y(N152) );
  MXI4X1 U2346 ( .A(\CACHE[4][35] ), .B(\CACHE[5][35] ), .C(\CACHE[6][35] ), 
        .D(\CACHE[7][35] ), .S0(n428), .S1(n450), .Y(n3167) );
  MXI4X1 U2347 ( .A(\CACHE[0][35] ), .B(\CACHE[1][35] ), .C(\CACHE[2][35] ), 
        .D(\CACHE[3][35] ), .S0(n428), .S1(n452), .Y(n3166) );
  MXI2X1 U2348 ( .A(n3168), .B(n3169), .S0(n465), .Y(N151) );
  MXI4X1 U2349 ( .A(\CACHE[4][36] ), .B(\CACHE[5][36] ), .C(\CACHE[6][36] ), 
        .D(\CACHE[7][36] ), .S0(n428), .S1(n443), .Y(n3169) );
  MXI4X1 U2350 ( .A(\CACHE[0][36] ), .B(\CACHE[1][36] ), .C(\CACHE[2][36] ), 
        .D(\CACHE[3][36] ), .S0(n428), .S1(n443), .Y(n3168) );
  MXI2X1 U2351 ( .A(n3170), .B(n3171), .S0(n465), .Y(N150) );
  MXI4X1 U2352 ( .A(\CACHE[4][37] ), .B(\CACHE[5][37] ), .C(\CACHE[6][37] ), 
        .D(\CACHE[7][37] ), .S0(n428), .S1(n443), .Y(n3171) );
  MXI4X1 U2353 ( .A(\CACHE[0][37] ), .B(\CACHE[1][37] ), .C(\CACHE[2][37] ), 
        .D(\CACHE[3][37] ), .S0(n428), .S1(n443), .Y(n3170) );
  MXI2X1 U2354 ( .A(n3172), .B(n3173), .S0(n465), .Y(N149) );
  MXI4X1 U2355 ( .A(\CACHE[4][38] ), .B(\CACHE[5][38] ), .C(\CACHE[6][38] ), 
        .D(\CACHE[7][38] ), .S0(n428), .S1(n443), .Y(n3173) );
  MXI4X1 U2356 ( .A(\CACHE[0][38] ), .B(\CACHE[1][38] ), .C(\CACHE[2][38] ), 
        .D(\CACHE[3][38] ), .S0(n428), .S1(n443), .Y(n3172) );
  MXI2X1 U2357 ( .A(n3174), .B(n3175), .S0(n465), .Y(N148) );
  MXI4X1 U2358 ( .A(\CACHE[4][39] ), .B(\CACHE[5][39] ), .C(\CACHE[6][39] ), 
        .D(\CACHE[7][39] ), .S0(n428), .S1(n443), .Y(n3175) );
  MXI4X1 U2359 ( .A(\CACHE[0][39] ), .B(\CACHE[1][39] ), .C(\CACHE[2][39] ), 
        .D(\CACHE[3][39] ), .S0(n429), .S1(n443), .Y(n3174) );
  MXI2X1 U2360 ( .A(n3176), .B(n3177), .S0(n465), .Y(N147) );
  MXI4X1 U2361 ( .A(\CACHE[4][40] ), .B(\CACHE[5][40] ), .C(\CACHE[6][40] ), 
        .D(\CACHE[7][40] ), .S0(n429), .S1(n443), .Y(n3177) );
  MXI4X1 U2362 ( .A(\CACHE[0][40] ), .B(\CACHE[1][40] ), .C(\CACHE[2][40] ), 
        .D(\CACHE[3][40] ), .S0(n429), .S1(n443), .Y(n3176) );
  MXI2X1 U2363 ( .A(n3178), .B(n3179), .S0(n465), .Y(N146) );
  MXI4X1 U2364 ( .A(\CACHE[4][41] ), .B(\CACHE[5][41] ), .C(\CACHE[6][41] ), 
        .D(\CACHE[7][41] ), .S0(n429), .S1(n443), .Y(n3179) );
  MXI4X1 U2365 ( .A(\CACHE[0][41] ), .B(\CACHE[1][41] ), .C(\CACHE[2][41] ), 
        .D(\CACHE[3][41] ), .S0(n429), .S1(n443), .Y(n3178) );
  MXI2X1 U2366 ( .A(n3180), .B(n3181), .S0(n465), .Y(N145) );
  MXI4X1 U2367 ( .A(\CACHE[4][42] ), .B(\CACHE[5][42] ), .C(\CACHE[6][42] ), 
        .D(\CACHE[7][42] ), .S0(n429), .S1(n450), .Y(n3181) );
  MXI4X1 U2368 ( .A(\CACHE[0][42] ), .B(\CACHE[1][42] ), .C(\CACHE[2][42] ), 
        .D(\CACHE[3][42] ), .S0(n429), .S1(n452), .Y(n3180) );
  MXI2X1 U2369 ( .A(n3182), .B(n3183), .S0(n465), .Y(N144) );
  MXI4X1 U2370 ( .A(\CACHE[4][43] ), .B(\CACHE[5][43] ), .C(\CACHE[6][43] ), 
        .D(\CACHE[7][43] ), .S0(n429), .S1(n448), .Y(n3183) );
  MXI4X1 U2371 ( .A(\CACHE[0][43] ), .B(\CACHE[1][43] ), .C(\CACHE[2][43] ), 
        .D(\CACHE[3][43] ), .S0(n429), .S1(n443), .Y(n3182) );
  MXI2X1 U2372 ( .A(n3184), .B(n3185), .S0(n465), .Y(N143) );
  MXI4X1 U2373 ( .A(\CACHE[4][44] ), .B(\CACHE[5][44] ), .C(\CACHE[6][44] ), 
        .D(\CACHE[7][44] ), .S0(n429), .S1(n444), .Y(n3185) );
  MXI4X1 U2374 ( .A(\CACHE[0][44] ), .B(\CACHE[1][44] ), .C(\CACHE[2][44] ), 
        .D(\CACHE[3][44] ), .S0(n429), .S1(n451), .Y(n3184) );
  MXI2X1 U2375 ( .A(n3186), .B(n3187), .S0(n465), .Y(N142) );
  MXI4X1 U2376 ( .A(\CACHE[4][45] ), .B(\CACHE[5][45] ), .C(\CACHE[6][45] ), 
        .D(\CACHE[7][45] ), .S0(n429), .S1(n455), .Y(n3187) );
  MXI4X1 U2377 ( .A(\CACHE[0][45] ), .B(\CACHE[1][45] ), .C(\CACHE[2][45] ), 
        .D(\CACHE[3][45] ), .S0(n429), .S1(n453), .Y(n3186) );
  MXI2X1 U2378 ( .A(n3188), .B(n3189), .S0(n465), .Y(N141) );
  MXI4X1 U2379 ( .A(\CACHE[4][46] ), .B(\CACHE[5][46] ), .C(\CACHE[6][46] ), 
        .D(\CACHE[7][46] ), .S0(n430), .S1(n457), .Y(n3189) );
  MXI4X1 U2380 ( .A(\CACHE[0][46] ), .B(\CACHE[1][46] ), .C(\CACHE[2][46] ), 
        .D(\CACHE[3][46] ), .S0(n430), .S1(n454), .Y(n3188) );
  MXI2X1 U2381 ( .A(n3190), .B(n3191), .S0(n465), .Y(N140) );
  MXI4X1 U2382 ( .A(\CACHE[4][47] ), .B(\CACHE[5][47] ), .C(\CACHE[6][47] ), 
        .D(\CACHE[7][47] ), .S0(n430), .S1(n442), .Y(n3191) );
  MXI4X1 U2383 ( .A(\CACHE[0][47] ), .B(\CACHE[1][47] ), .C(\CACHE[2][47] ), 
        .D(\CACHE[3][47] ), .S0(n430), .S1(n441), .Y(n3190) );
  MXI2X1 U2384 ( .A(n3192), .B(n3193), .S0(n463), .Y(N139) );
  MXI4X1 U2385 ( .A(\CACHE[4][48] ), .B(\CACHE[5][48] ), .C(\CACHE[6][48] ), 
        .D(\CACHE[7][48] ), .S0(n430), .S1(n444), .Y(n3193) );
  MXI4X1 U2386 ( .A(\CACHE[0][48] ), .B(\CACHE[1][48] ), .C(\CACHE[2][48] ), 
        .D(\CACHE[3][48] ), .S0(n430), .S1(n444), .Y(n3192) );
  MXI2X1 U2387 ( .A(n3194), .B(n3195), .S0(n464), .Y(N138) );
  MXI4X1 U2388 ( .A(\CACHE[4][49] ), .B(\CACHE[5][49] ), .C(\CACHE[6][49] ), 
        .D(\CACHE[7][49] ), .S0(n430), .S1(n444), .Y(n3195) );
  MXI4X1 U2389 ( .A(\CACHE[0][49] ), .B(\CACHE[1][49] ), .C(\CACHE[2][49] ), 
        .D(\CACHE[3][49] ), .S0(n430), .S1(n444), .Y(n3194) );
  MXI2X1 U2390 ( .A(n3196), .B(n3197), .S0(n466), .Y(N137) );
  MXI4X1 U2391 ( .A(\CACHE[4][50] ), .B(\CACHE[5][50] ), .C(\CACHE[6][50] ), 
        .D(\CACHE[7][50] ), .S0(n430), .S1(n444), .Y(n3197) );
  MXI4X1 U2392 ( .A(\CACHE[0][50] ), .B(\CACHE[1][50] ), .C(\CACHE[2][50] ), 
        .D(\CACHE[3][50] ), .S0(n430), .S1(n444), .Y(n3196) );
  MXI2X1 U2393 ( .A(n3198), .B(n3199), .S0(n467), .Y(N136) );
  MXI4X1 U2394 ( .A(\CACHE[4][51] ), .B(\CACHE[5][51] ), .C(\CACHE[6][51] ), 
        .D(\CACHE[7][51] ), .S0(n430), .S1(n444), .Y(n3199) );
  MXI4X1 U2395 ( .A(\CACHE[0][51] ), .B(\CACHE[1][51] ), .C(\CACHE[2][51] ), 
        .D(\CACHE[3][51] ), .S0(n430), .S1(n444), .Y(n3198) );
  MXI2X1 U2396 ( .A(n3200), .B(n3201), .S0(n468), .Y(N135) );
  MXI4X1 U2397 ( .A(\CACHE[4][52] ), .B(\CACHE[5][52] ), .C(\CACHE[6][52] ), 
        .D(\CACHE[7][52] ), .S0(n431), .S1(n444), .Y(n3201) );
  MXI4X1 U2398 ( .A(\CACHE[0][52] ), .B(\CACHE[1][52] ), .C(\CACHE[2][52] ), 
        .D(\CACHE[3][52] ), .S0(n431), .S1(n444), .Y(n3200) );
  MXI2X1 U2399 ( .A(n3202), .B(n3203), .S0(n465), .Y(N134) );
  MXI4X1 U2400 ( .A(\CACHE[4][53] ), .B(\CACHE[5][53] ), .C(\CACHE[6][53] ), 
        .D(\CACHE[7][53] ), .S0(n430), .S1(n444), .Y(n3203) );
  MXI4X1 U2401 ( .A(\CACHE[0][53] ), .B(\CACHE[1][53] ), .C(\CACHE[2][53] ), 
        .D(\CACHE[3][53] ), .S0(n431), .S1(n444), .Y(n3202) );
  MXI2X1 U2402 ( .A(n3204), .B(n3205), .S0(n470), .Y(N133) );
  MXI4X1 U2403 ( .A(\CACHE[4][54] ), .B(\CACHE[5][54] ), .C(\CACHE[6][54] ), 
        .D(\CACHE[7][54] ), .S0(n431), .S1(n445), .Y(n3205) );
  MXI4X1 U2404 ( .A(\CACHE[0][54] ), .B(\CACHE[1][54] ), .C(\CACHE[2][54] ), 
        .D(\CACHE[3][54] ), .S0(n431), .S1(n445), .Y(n3204) );
  MXI2X1 U2405 ( .A(n3206), .B(n3207), .S0(n469), .Y(N132) );
  MXI4X1 U2406 ( .A(\CACHE[4][55] ), .B(\CACHE[5][55] ), .C(\CACHE[6][55] ), 
        .D(\CACHE[7][55] ), .S0(n431), .S1(n445), .Y(n3207) );
  MXI4X1 U2407 ( .A(\CACHE[0][55] ), .B(\CACHE[1][55] ), .C(\CACHE[2][55] ), 
        .D(\CACHE[3][55] ), .S0(n431), .S1(n445), .Y(n3206) );
  MXI2X1 U2408 ( .A(n3208), .B(n3209), .S0(n462), .Y(N131) );
  MXI4X1 U2409 ( .A(\CACHE[4][56] ), .B(\CACHE[5][56] ), .C(\CACHE[6][56] ), 
        .D(\CACHE[7][56] ), .S0(n431), .S1(n445), .Y(n3209) );
  MXI4X1 U2410 ( .A(\CACHE[0][56] ), .B(\CACHE[1][56] ), .C(\CACHE[2][56] ), 
        .D(\CACHE[3][56] ), .S0(n431), .S1(n445), .Y(n3208) );
  MXI2X1 U2411 ( .A(n3210), .B(n3211), .S0(n463), .Y(N130) );
  MXI4X1 U2412 ( .A(\CACHE[4][57] ), .B(\CACHE[5][57] ), .C(\CACHE[6][57] ), 
        .D(\CACHE[7][57] ), .S0(n431), .S1(n445), .Y(n3211) );
  MXI4X1 U2413 ( .A(\CACHE[0][57] ), .B(\CACHE[1][57] ), .C(\CACHE[2][57] ), 
        .D(\CACHE[3][57] ), .S0(n431), .S1(n445), .Y(n3210) );
  MXI2X1 U2414 ( .A(n3212), .B(n3213), .S0(n464), .Y(N129) );
  MXI4X1 U2415 ( .A(\CACHE[4][58] ), .B(\CACHE[5][58] ), .C(\CACHE[6][58] ), 
        .D(\CACHE[7][58] ), .S0(n431), .S1(n445), .Y(n3213) );
  MXI4X1 U2416 ( .A(\CACHE[0][58] ), .B(\CACHE[1][58] ), .C(\CACHE[2][58] ), 
        .D(\CACHE[3][58] ), .S0(n432), .S1(n445), .Y(n3212) );
  MXI2X1 U2417 ( .A(n3214), .B(n3215), .S0(n466), .Y(N128) );
  MXI4X1 U2418 ( .A(\CACHE[4][59] ), .B(\CACHE[5][59] ), .C(\CACHE[6][59] ), 
        .D(\CACHE[7][59] ), .S0(n431), .S1(n445), .Y(n3215) );
  MXI4X1 U2419 ( .A(\CACHE[0][59] ), .B(\CACHE[1][59] ), .C(\CACHE[2][59] ), 
        .D(\CACHE[3][59] ), .S0(n432), .S1(n445), .Y(n3214) );
  MXI2X1 U2420 ( .A(n3216), .B(n3217), .S0(n465), .Y(N127) );
  MXI4X1 U2421 ( .A(\CACHE[4][60] ), .B(\CACHE[5][60] ), .C(\CACHE[6][60] ), 
        .D(\CACHE[7][60] ), .S0(n432), .S1(n446), .Y(n3217) );
  MXI4X1 U2422 ( .A(\CACHE[0][60] ), .B(\CACHE[1][60] ), .C(\CACHE[2][60] ), 
        .D(\CACHE[3][60] ), .S0(n432), .S1(n446), .Y(n3216) );
  MXI2X1 U2423 ( .A(n3218), .B(n3219), .S0(n470), .Y(N126) );
  MXI4X1 U2424 ( .A(\CACHE[4][61] ), .B(\CACHE[5][61] ), .C(\CACHE[6][61] ), 
        .D(\CACHE[7][61] ), .S0(n432), .S1(n446), .Y(n3219) );
  MXI4X1 U2425 ( .A(\CACHE[0][61] ), .B(\CACHE[1][61] ), .C(\CACHE[2][61] ), 
        .D(\CACHE[3][61] ), .S0(n432), .S1(n446), .Y(n3218) );
  MXI2X1 U2426 ( .A(n3220), .B(n3221), .S0(n470), .Y(N125) );
  MXI4X1 U2427 ( .A(\CACHE[4][62] ), .B(\CACHE[5][62] ), .C(\CACHE[6][62] ), 
        .D(\CACHE[7][62] ), .S0(n432), .S1(n446), .Y(n3221) );
  MXI4X1 U2428 ( .A(\CACHE[0][62] ), .B(\CACHE[1][62] ), .C(\CACHE[2][62] ), 
        .D(\CACHE[3][62] ), .S0(n432), .S1(n446), .Y(n3220) );
  MXI2X1 U2429 ( .A(n3222), .B(n3223), .S0(n469), .Y(N124) );
  MXI4X1 U2430 ( .A(\CACHE[4][63] ), .B(\CACHE[5][63] ), .C(\CACHE[6][63] ), 
        .D(\CACHE[7][63] ), .S0(n432), .S1(n446), .Y(n3223) );
  MXI4X1 U2431 ( .A(\CACHE[0][63] ), .B(\CACHE[1][63] ), .C(\CACHE[2][63] ), 
        .D(\CACHE[3][63] ), .S0(n432), .S1(n446), .Y(n3222) );
  MXI2X1 U2432 ( .A(n3224), .B(n3225), .S0(n462), .Y(N123) );
  MXI4X1 U2433 ( .A(\CACHE[4][64] ), .B(\CACHE[5][64] ), .C(\CACHE[6][64] ), 
        .D(\CACHE[7][64] ), .S0(n432), .S1(n446), .Y(n3225) );
  MXI4X1 U2434 ( .A(\CACHE[0][64] ), .B(\CACHE[1][64] ), .C(\CACHE[2][64] ), 
        .D(\CACHE[3][64] ), .S0(n432), .S1(n446), .Y(n3224) );
  MXI2X1 U2435 ( .A(n3226), .B(n3227), .S0(n463), .Y(N122) );
  MXI4X1 U2436 ( .A(\CACHE[4][65] ), .B(\CACHE[5][65] ), .C(\CACHE[6][65] ), 
        .D(\CACHE[7][65] ), .S0(n432), .S1(n446), .Y(n3227) );
  MXI4X1 U2437 ( .A(\CACHE[0][65] ), .B(\CACHE[1][65] ), .C(\CACHE[2][65] ), 
        .D(\CACHE[3][65] ), .S0(n433), .S1(n446), .Y(n3226) );
  MXI2X1 U2438 ( .A(n3228), .B(n3229), .S0(n464), .Y(N121) );
  MXI4X1 U2439 ( .A(\CACHE[4][66] ), .B(\CACHE[5][66] ), .C(\CACHE[6][66] ), 
        .D(\CACHE[7][66] ), .S0(n433), .S1(n447), .Y(n3229) );
  MXI4X1 U2440 ( .A(\CACHE[0][66] ), .B(\CACHE[1][66] ), .C(\CACHE[2][66] ), 
        .D(\CACHE[3][66] ), .S0(n433), .S1(n447), .Y(n3228) );
  MXI2X1 U2441 ( .A(n3230), .B(n3231), .S0(n466), .Y(N120) );
  MXI4X1 U2442 ( .A(\CACHE[4][67] ), .B(\CACHE[5][67] ), .C(\CACHE[6][67] ), 
        .D(\CACHE[7][67] ), .S0(n433), .S1(n447), .Y(n3231) );
  MXI4X1 U2443 ( .A(\CACHE[0][67] ), .B(\CACHE[1][67] ), .C(\CACHE[2][67] ), 
        .D(\CACHE[3][67] ), .S0(n433), .S1(n447), .Y(n3230) );
  MXI2X1 U2444 ( .A(n3232), .B(n3233), .S0(n467), .Y(N119) );
  MXI4X1 U2445 ( .A(\CACHE[4][68] ), .B(\CACHE[5][68] ), .C(\CACHE[6][68] ), 
        .D(\CACHE[7][68] ), .S0(n433), .S1(n447), .Y(n3233) );
  MXI4X1 U2446 ( .A(\CACHE[0][68] ), .B(\CACHE[1][68] ), .C(\CACHE[2][68] ), 
        .D(\CACHE[3][68] ), .S0(n433), .S1(n447), .Y(n3232) );
  MXI2X1 U2447 ( .A(n3234), .B(n3235), .S0(n468), .Y(N118) );
  MXI4X1 U2448 ( .A(\CACHE[4][69] ), .B(\CACHE[5][69] ), .C(\CACHE[6][69] ), 
        .D(\CACHE[7][69] ), .S0(n433), .S1(n447), .Y(n3235) );
  MXI4X1 U2449 ( .A(\CACHE[0][69] ), .B(\CACHE[1][69] ), .C(\CACHE[2][69] ), 
        .D(\CACHE[3][69] ), .S0(n433), .S1(n447), .Y(n3234) );
  MXI2X1 U2450 ( .A(n3236), .B(n3237), .S0(n465), .Y(N117) );
  MXI4X1 U2451 ( .A(\CACHE[4][70] ), .B(\CACHE[5][70] ), .C(\CACHE[6][70] ), 
        .D(\CACHE[7][70] ), .S0(n433), .S1(n447), .Y(n3237) );
  MXI4X1 U2452 ( .A(\CACHE[0][70] ), .B(\CACHE[1][70] ), .C(\CACHE[2][70] ), 
        .D(\CACHE[3][70] ), .S0(n433), .S1(n447), .Y(n3236) );
  MXI2X1 U2453 ( .A(n3238), .B(n3239), .S0(n469), .Y(N116) );
  MXI4X1 U2454 ( .A(\CACHE[4][71] ), .B(\CACHE[5][71] ), .C(\CACHE[6][71] ), 
        .D(\CACHE[7][71] ), .S0(n433), .S1(n447), .Y(n3239) );
  MXI4X1 U2455 ( .A(\CACHE[0][71] ), .B(\CACHE[1][71] ), .C(\CACHE[2][71] ), 
        .D(\CACHE[3][71] ), .S0(n434), .S1(n447), .Y(n3238) );
  MXI2X1 U2456 ( .A(n3240), .B(n3241), .S0(n467), .Y(N115) );
  MXI4X1 U2457 ( .A(\CACHE[4][72] ), .B(\CACHE[5][72] ), .C(\CACHE[6][72] ), 
        .D(\CACHE[7][72] ), .S0(n434), .S1(n445), .Y(n3241) );
  MXI4X1 U2458 ( .A(\CACHE[0][72] ), .B(\CACHE[1][72] ), .C(\CACHE[2][72] ), 
        .D(\CACHE[3][72] ), .S0(n433), .S1(n449), .Y(n3240) );
  MXI2X1 U2459 ( .A(n3242), .B(n3243), .S0(n468), .Y(N114) );
  MXI4X1 U2460 ( .A(\CACHE[4][73] ), .B(\CACHE[5][73] ), .C(\CACHE[6][73] ), 
        .D(\CACHE[7][73] ), .S0(n434), .S1(n447), .Y(n3243) );
  MXI4X1 U2461 ( .A(\CACHE[0][73] ), .B(\CACHE[1][73] ), .C(\CACHE[2][73] ), 
        .D(\CACHE[3][73] ), .S0(n434), .S1(n446), .Y(n3242) );
  MXI2X1 U2462 ( .A(n3244), .B(n3245), .S0(n465), .Y(N113) );
  MXI4X1 U2463 ( .A(\CACHE[4][74] ), .B(\CACHE[5][74] ), .C(\CACHE[6][74] ), 
        .D(\CACHE[7][74] ), .S0(n434), .S1(n439), .Y(n3245) );
  MXI4X1 U2464 ( .A(\CACHE[0][74] ), .B(\CACHE[1][74] ), .C(\CACHE[2][74] ), 
        .D(\CACHE[3][74] ), .S0(n434), .S1(n456), .Y(n3244) );
  MXI2X1 U2465 ( .A(n3246), .B(n3247), .S0(n462), .Y(N112) );
  MXI4X1 U2466 ( .A(\CACHE[4][75] ), .B(\CACHE[5][75] ), .C(\CACHE[6][75] ), 
        .D(\CACHE[7][75] ), .S0(n434), .S1(n453), .Y(n3247) );
  MXI4X1 U2467 ( .A(\CACHE[0][75] ), .B(\CACHE[1][75] ), .C(\CACHE[2][75] ), 
        .D(\CACHE[3][75] ), .S0(n434), .S1(n444), .Y(n3246) );
  MXI2X1 U2468 ( .A(n3248), .B(n3249), .S0(n468), .Y(N111) );
  MXI4X1 U2469 ( .A(\CACHE[4][76] ), .B(\CACHE[5][76] ), .C(\CACHE[6][76] ), 
        .D(\CACHE[7][76] ), .S0(n434), .S1(n457), .Y(n3249) );
  MXI4X1 U2470 ( .A(\CACHE[0][76] ), .B(\CACHE[1][76] ), .C(\CACHE[2][76] ), 
        .D(\CACHE[3][76] ), .S0(n434), .S1(n455), .Y(n3248) );
  MXI2X1 U2471 ( .A(n3250), .B(n3251), .S0(n470), .Y(N110) );
  MXI4X1 U2472 ( .A(\CACHE[4][77] ), .B(\CACHE[5][77] ), .C(\CACHE[6][77] ), 
        .D(\CACHE[7][77] ), .S0(n434), .S1(n442), .Y(n3251) );
  MXI4X1 U2473 ( .A(\CACHE[0][77] ), .B(\CACHE[1][77] ), .C(\CACHE[2][77] ), 
        .D(\CACHE[3][77] ), .S0(n434), .S1(n441), .Y(n3250) );
  MXI2X1 U2474 ( .A(n3252), .B(n3253), .S0(n469), .Y(N109) );
  MXI4X1 U2475 ( .A(\CACHE[4][78] ), .B(\CACHE[5][78] ), .C(\CACHE[6][78] ), 
        .D(\CACHE[7][78] ), .S0(n415), .S1(n448), .Y(n3253) );
  MXI4X1 U2476 ( .A(\CACHE[0][78] ), .B(\CACHE[1][78] ), .C(\CACHE[2][78] ), 
        .D(\CACHE[3][78] ), .S0(n415), .S1(n448), .Y(n3252) );
  MXI2X1 U2477 ( .A(n3254), .B(n3255), .S0(n462), .Y(N108) );
  MXI4X1 U2478 ( .A(\CACHE[4][79] ), .B(\CACHE[5][79] ), .C(\CACHE[6][79] ), 
        .D(\CACHE[7][79] ), .S0(n415), .S1(n448), .Y(n3255) );
  MXI4X1 U2479 ( .A(\CACHE[0][79] ), .B(\CACHE[1][79] ), .C(\CACHE[2][79] ), 
        .D(\CACHE[3][79] ), .S0(n415), .S1(n448), .Y(n3254) );
  MXI2X1 U2480 ( .A(n3256), .B(n3257), .S0(n463), .Y(N107) );
  MXI4X1 U2481 ( .A(\CACHE[4][80] ), .B(\CACHE[5][80] ), .C(\CACHE[6][80] ), 
        .D(\CACHE[7][80] ), .S0(n415), .S1(n448), .Y(n3257) );
  MXI4X1 U2482 ( .A(\CACHE[0][80] ), .B(\CACHE[1][80] ), .C(\CACHE[2][80] ), 
        .D(\CACHE[3][80] ), .S0(n415), .S1(n448), .Y(n3256) );
  MXI2X1 U2483 ( .A(n3258), .B(n3259), .S0(n464), .Y(N106) );
  MXI4X1 U2484 ( .A(\CACHE[4][81] ), .B(\CACHE[5][81] ), .C(\CACHE[6][81] ), 
        .D(\CACHE[7][81] ), .S0(n415), .S1(n448), .Y(n3259) );
  MXI4X1 U2485 ( .A(\CACHE[0][81] ), .B(\CACHE[1][81] ), .C(\CACHE[2][81] ), 
        .D(\CACHE[3][81] ), .S0(n415), .S1(n448), .Y(n3258) );
  MXI2X1 U2486 ( .A(n3260), .B(n3261), .S0(n466), .Y(N105) );
  MXI4X1 U2487 ( .A(\CACHE[4][82] ), .B(\CACHE[5][82] ), .C(\CACHE[6][82] ), 
        .D(\CACHE[7][82] ), .S0(n415), .S1(n448), .Y(n3261) );
  MXI4X1 U2488 ( .A(\CACHE[0][82] ), .B(\CACHE[1][82] ), .C(\CACHE[2][82] ), 
        .D(\CACHE[3][82] ), .S0(n415), .S1(n448), .Y(n3260) );
  MXI2X1 U2489 ( .A(n3262), .B(n3263), .S0(n467), .Y(N104) );
  MXI4X1 U2490 ( .A(\CACHE[4][83] ), .B(\CACHE[5][83] ), .C(\CACHE[6][83] ), 
        .D(\CACHE[7][83] ), .S0(n415), .S1(n448), .Y(n3263) );
  MXI4X1 U2491 ( .A(\CACHE[0][83] ), .B(\CACHE[1][83] ), .C(\CACHE[2][83] ), 
        .D(\CACHE[3][83] ), .S0(n415), .S1(n448), .Y(n3262) );
  MXI2X1 U2492 ( .A(n3264), .B(n3265), .S0(n471), .Y(N103) );
  MXI4X1 U2493 ( .A(\CACHE[4][84] ), .B(\CACHE[5][84] ), .C(\CACHE[6][84] ), 
        .D(\CACHE[7][84] ), .S0(n416), .S1(n449), .Y(n3265) );
  MXI4X1 U2494 ( .A(\CACHE[0][84] ), .B(\CACHE[1][84] ), .C(\CACHE[2][84] ), 
        .D(\CACHE[3][84] ), .S0(n416), .S1(n449), .Y(n3264) );
  MXI2X1 U2495 ( .A(n3266), .B(n3267), .S0(N32), .Y(N102) );
  MXI4X1 U2496 ( .A(\CACHE[4][85] ), .B(\CACHE[5][85] ), .C(\CACHE[6][85] ), 
        .D(\CACHE[7][85] ), .S0(n416), .S1(n449), .Y(n3267) );
  MXI4X1 U2497 ( .A(\CACHE[0][85] ), .B(\CACHE[1][85] ), .C(\CACHE[2][85] ), 
        .D(\CACHE[3][85] ), .S0(n416), .S1(n449), .Y(n3266) );
  MXI2X1 U2498 ( .A(n3268), .B(n3269), .S0(n471), .Y(N101) );
  MXI4X1 U2499 ( .A(\CACHE[4][86] ), .B(\CACHE[5][86] ), .C(\CACHE[6][86] ), 
        .D(\CACHE[7][86] ), .S0(n416), .S1(n449), .Y(n3269) );
  MXI4X1 U2500 ( .A(\CACHE[0][86] ), .B(\CACHE[1][86] ), .C(\CACHE[2][86] ), 
        .D(\CACHE[3][86] ), .S0(n416), .S1(n449), .Y(n3268) );
  MXI2X1 U2501 ( .A(n3270), .B(n3271), .S0(N32), .Y(N100) );
  MXI4X1 U2502 ( .A(\CACHE[4][87] ), .B(\CACHE[5][87] ), .C(\CACHE[6][87] ), 
        .D(\CACHE[7][87] ), .S0(n416), .S1(n449), .Y(n3271) );
  MXI4X1 U2503 ( .A(\CACHE[0][87] ), .B(\CACHE[1][87] ), .C(\CACHE[2][87] ), 
        .D(\CACHE[3][87] ), .S0(n416), .S1(n449), .Y(n3270) );
  MXI2X1 U2504 ( .A(n3272), .B(n3273), .S0(n471), .Y(N99) );
  MXI4X1 U2505 ( .A(\CACHE[4][88] ), .B(\CACHE[5][88] ), .C(\CACHE[6][88] ), 
        .D(\CACHE[7][88] ), .S0(n416), .S1(n449), .Y(n3273) );
  MXI4X1 U2506 ( .A(\CACHE[0][88] ), .B(\CACHE[1][88] ), .C(\CACHE[2][88] ), 
        .D(\CACHE[3][88] ), .S0(n416), .S1(n449), .Y(n3272) );
  MXI2X1 U2507 ( .A(n3274), .B(n3275), .S0(N32), .Y(N98) );
  MXI4X1 U2508 ( .A(\CACHE[4][89] ), .B(\CACHE[5][89] ), .C(\CACHE[6][89] ), 
        .D(\CACHE[7][89] ), .S0(n416), .S1(n449), .Y(n3275) );
  MXI4X1 U2509 ( .A(\CACHE[0][89] ), .B(\CACHE[1][89] ), .C(\CACHE[2][89] ), 
        .D(\CACHE[3][89] ), .S0(n416), .S1(n449), .Y(n3274) );
  MXI2X1 U2510 ( .A(n3276), .B(n3277), .S0(n471), .Y(N97) );
  MXI4X1 U2511 ( .A(\CACHE[4][90] ), .B(\CACHE[5][90] ), .C(\CACHE[6][90] ), 
        .D(\CACHE[7][90] ), .S0(n416), .S1(n450), .Y(n3277) );
  MXI4X1 U2512 ( .A(\CACHE[0][90] ), .B(\CACHE[1][90] ), .C(\CACHE[2][90] ), 
        .D(\CACHE[3][90] ), .S0(n426), .S1(n450), .Y(n3276) );
  MXI2X1 U2513 ( .A(n3278), .B(n3279), .S0(n469), .Y(N96) );
  MXI4X1 U2514 ( .A(\CACHE[4][91] ), .B(\CACHE[5][91] ), .C(\CACHE[6][91] ), 
        .D(\CACHE[7][91] ), .S0(n430), .S1(n450), .Y(n3279) );
  MXI4X1 U2515 ( .A(\CACHE[0][91] ), .B(\CACHE[1][91] ), .C(\CACHE[2][91] ), 
        .D(\CACHE[3][91] ), .S0(n434), .S1(n450), .Y(n3278) );
  MXI2X1 U2516 ( .A(n3280), .B(n3281), .S0(n462), .Y(N95) );
  MXI4X1 U2517 ( .A(\CACHE[4][92] ), .B(\CACHE[5][92] ), .C(\CACHE[6][92] ), 
        .D(\CACHE[7][92] ), .S0(n423), .S1(n450), .Y(n3281) );
  MXI4X1 U2518 ( .A(\CACHE[0][92] ), .B(\CACHE[1][92] ), .C(\CACHE[2][92] ), 
        .D(\CACHE[3][92] ), .S0(n431), .S1(n450), .Y(n3280) );
  MXI2X1 U2519 ( .A(n3282), .B(n3283), .S0(n463), .Y(N94) );
  MXI4X1 U2520 ( .A(\CACHE[4][93] ), .B(\CACHE[5][93] ), .C(\CACHE[6][93] ), 
        .D(\CACHE[7][93] ), .S0(n421), .S1(n450), .Y(n3283) );
  MXI4X1 U2521 ( .A(\CACHE[0][93] ), .B(\CACHE[1][93] ), .C(\CACHE[2][93] ), 
        .D(\CACHE[3][93] ), .S0(n426), .S1(n450), .Y(n3282) );
  MXI2X1 U2522 ( .A(n3284), .B(n3285), .S0(n464), .Y(N93) );
  MXI4X1 U2523 ( .A(\CACHE[4][94] ), .B(\CACHE[5][94] ), .C(\CACHE[6][94] ), 
        .D(\CACHE[7][94] ), .S0(n433), .S1(n450), .Y(n3285) );
  MXI4X1 U2524 ( .A(\CACHE[0][94] ), .B(\CACHE[1][94] ), .C(\CACHE[2][94] ), 
        .D(\CACHE[3][94] ), .S0(n422), .S1(n450), .Y(n3284) );
  MXI2X1 U2525 ( .A(n3286), .B(n3287), .S0(n466), .Y(N92) );
  MXI4X1 U2526 ( .A(\CACHE[4][95] ), .B(\CACHE[5][95] ), .C(\CACHE[6][95] ), 
        .D(\CACHE[7][95] ), .S0(n424), .S1(n450), .Y(n3287) );
  MXI4X1 U2527 ( .A(\CACHE[0][95] ), .B(\CACHE[1][95] ), .C(\CACHE[2][95] ), 
        .D(\CACHE[3][95] ), .S0(n425), .S1(n450), .Y(n3286) );
  NAND3BX1 U2528 ( .AN(n3404), .B(n3405), .C(n3406), .Y(proc_stall) );
  OAI221XL U2529 ( .A0(n3407), .A1(n3408), .B0(n3409), .B1(n3410), .C0(n3411), 
        .Y(proc_rdata[9]) );
  OAI221XL U2530 ( .A0(n3407), .A1(n3416), .B0(n3409), .B1(n3417), .C0(n3418), 
        .Y(proc_rdata[8]) );
  OAI221XL U2531 ( .A0(n3407), .A1(n3421), .B0(n3409), .B1(n3422), .C0(n3423), 
        .Y(proc_rdata[7]) );
  OAI221XL U2532 ( .A0(n3407), .A1(n3426), .B0(n3409), .B1(n3427), .C0(n3428), 
        .Y(proc_rdata[6]) );
  OAI221XL U2533 ( .A0(n3407), .A1(n3431), .B0(n3409), .B1(n3432), .C0(n3433), 
        .Y(proc_rdata[5]) );
  OAI221XL U2534 ( .A0(n3407), .A1(n3436), .B0(n3409), .B1(n3437), .C0(n3438), 
        .Y(proc_rdata[4]) );
  OAI221XL U2535 ( .A0(n3407), .A1(n3441), .B0(n3409), .B1(n3442), .C0(n3443), 
        .Y(proc_rdata[3]) );
  OAI221XL U2536 ( .A0(n3407), .A1(n3446), .B0(n3409), .B1(n3447), .C0(n3448), 
        .Y(proc_rdata[31]) );
  OAI221XL U2537 ( .A0(n3407), .A1(n3451), .B0(n3409), .B1(n3452), .C0(n3453), 
        .Y(proc_rdata[30]) );
  OAI221XL U2538 ( .A0(n3407), .A1(n3456), .B0(n3409), .B1(n3457), .C0(n3458), 
        .Y(proc_rdata[2]) );
  OAI221XL U2539 ( .A0(n3407), .A1(n3461), .B0(n3409), .B1(n3462), .C0(n3463), 
        .Y(proc_rdata[29]) );
  OAI221XL U2540 ( .A0(n3407), .A1(n3466), .B0(n3409), .B1(n3467), .C0(n3468), 
        .Y(proc_rdata[28]) );
  OAI221XL U2541 ( .A0(n3407), .A1(n3471), .B0(n3409), .B1(n3472), .C0(n3473), 
        .Y(proc_rdata[27]) );
  OAI221XL U2542 ( .A0(n3407), .A1(n3476), .B0(n3409), .B1(n3477), .C0(n3478), 
        .Y(proc_rdata[26]) );
  OAI221XL U2543 ( .A0(n3407), .A1(n3481), .B0(n3409), .B1(n3482), .C0(n3483), 
        .Y(proc_rdata[25]) );
  OAI221XL U2544 ( .A0(n3407), .A1(n3486), .B0(n3409), .B1(n3487), .C0(n3488), 
        .Y(proc_rdata[24]) );
  OAI221XL U2545 ( .A0(n3407), .A1(n3491), .B0(n3409), .B1(n3492), .C0(n3493), 
        .Y(proc_rdata[23]) );
  OAI221XL U2546 ( .A0(n3407), .A1(n3496), .B0(n3409), .B1(n3497), .C0(n3498), 
        .Y(proc_rdata[22]) );
  OAI221XL U2547 ( .A0(n3407), .A1(n3501), .B0(n3409), .B1(n3502), .C0(n3503), 
        .Y(proc_rdata[21]) );
  OAI221XL U2548 ( .A0(n3407), .A1(n3506), .B0(n3409), .B1(n3507), .C0(n3508), 
        .Y(proc_rdata[20]) );
  OAI221XL U2549 ( .A0(n3407), .A1(n3511), .B0(n3409), .B1(n3512), .C0(n3513), 
        .Y(proc_rdata[1]) );
  OAI221XL U2550 ( .A0(n3407), .A1(n3516), .B0(n3409), .B1(n3517), .C0(n3518), 
        .Y(proc_rdata[19]) );
  OAI221XL U2551 ( .A0(n3407), .A1(n3521), .B0(n3409), .B1(n3522), .C0(n3523), 
        .Y(proc_rdata[18]) );
  OAI221XL U2552 ( .A0(n3407), .A1(n3526), .B0(n3409), .B1(n3527), .C0(n3528), 
        .Y(proc_rdata[17]) );
  OAI221XL U2553 ( .A0(n3407), .A1(n3531), .B0(n3409), .B1(n3532), .C0(n3533), 
        .Y(proc_rdata[16]) );
  OAI221XL U2554 ( .A0(n3407), .A1(n3536), .B0(n3409), .B1(n3537), .C0(n3538), 
        .Y(proc_rdata[15]) );
  OAI221XL U2555 ( .A0(n3407), .A1(n3541), .B0(n3409), .B1(n3542), .C0(n3543), 
        .Y(proc_rdata[14]) );
  OAI221XL U2556 ( .A0(n3407), .A1(n3546), .B0(n3409), .B1(n3547), .C0(n3548), 
        .Y(proc_rdata[13]) );
  OAI221XL U2557 ( .A0(n3407), .A1(n3551), .B0(n3409), .B1(n3552), .C0(n3553), 
        .Y(proc_rdata[12]) );
  OAI221XL U2558 ( .A0(n3407), .A1(n3556), .B0(n3409), .B1(n3557), .C0(n3558), 
        .Y(proc_rdata[11]) );
  OAI221XL U2559 ( .A0(n3407), .A1(n3561), .B0(n3409), .B1(n3562), .C0(n3563), 
        .Y(proc_rdata[10]) );
  OAI221XL U2560 ( .A0(n3407), .A1(n3566), .B0(n3409), .B1(n3567), .C0(n3568), 
        .Y(proc_rdata[0]) );
  NOR3X1 U2561 ( .A(n460), .B(n435), .C(n472), .Y(n3575) );
  NOR3X1 U2562 ( .A(n460), .B(n434), .C(n472), .Y(n3730) );
  NOR3X1 U2563 ( .A(n436), .B(n458), .C(n472), .Y(n3731) );
  NOR3X1 U2564 ( .A(n422), .B(n458), .C(n472), .Y(n3732) );
  NOR3X1 U2565 ( .A(n435), .B(n470), .C(n459), .Y(n3733) );
  NOR3X1 U2566 ( .A(n421), .B(n470), .C(n459), .Y(n3734) );
  NOR3X1 U2567 ( .A(n458), .B(n471), .C(n437), .Y(n3735) );
  OAI31XL U2568 ( .A0(n3740), .A1(n3404), .A2(n3571), .B0(N34), .Y(n3738) );
  OAI31XL U2569 ( .A0(n3748), .A1(n3572), .A2(n3573), .B0(n3749), .Y(n3747) );
  OAI31XL U2570 ( .A0(n3748), .A1(proc_addr[0]), .A2(n3573), .B0(n3749), .Y(
        n3752) );
  OAI31XL U2571 ( .A0(n3748), .A1(proc_addr[1]), .A2(n3572), .B0(n3749), .Y(
        n3755) );
  NOR3X1 U2572 ( .A(n442), .B(n471), .C(n434), .Y(n3736) );
  OAI31XL U2573 ( .A0(n3748), .A1(proc_addr[1]), .A2(proc_addr[0]), .B0(n3749), 
        .Y(n3758) );
  NAND2BX1 U2574 ( .AN(n3748), .B(n3739), .Y(n3749) );
  NOR2X1 U2575 ( .A(n3759), .B(n3760), .Y(n3737) );
  CLKINVX1 U2576 ( .A(n3763), .Y(n3762) );
  AOI21X1 U2577 ( .A0(n3761), .A1(N34), .B0(n3740), .Y(n3743) );
  OAI31XL U2578 ( .A0(n3406), .A1(N34), .A2(n3404), .B0(n3405), .Y(n3764) );
  CLKINVX1 U2579 ( .A(N178), .Y(n3413) );
  CLKINVX1 U2580 ( .A(N88), .Y(n3445) );
  CLKINVX1 U2581 ( .A(N89), .Y(n3460) );
  CLKINVX1 U2582 ( .A(N90), .Y(n3515) );
  CLKINVX1 U2583 ( .A(N91), .Y(n3570) );
  CLKINVX1 U2584 ( .A(N92), .Y(n3446) );
  CLKINVX1 U2585 ( .A(N93), .Y(n3451) );
  CLKINVX1 U2586 ( .A(N94), .Y(n3461) );
  CLKINVX1 U2587 ( .A(N95), .Y(n3466) );
  CLKINVX1 U2588 ( .A(N96), .Y(n3471) );
  CLKINVX1 U2589 ( .A(N97), .Y(n3476) );
  CLKINVX1 U2590 ( .A(N179), .Y(n3419) );
  CLKINVX1 U2591 ( .A(N98), .Y(n3481) );
  CLKINVX1 U2592 ( .A(N99), .Y(n3486) );
  CLKINVX1 U2593 ( .A(N100), .Y(n3491) );
  CLKINVX1 U2594 ( .A(N101), .Y(n3496) );
  CLKINVX1 U2595 ( .A(N102), .Y(n3501) );
  CLKINVX1 U2596 ( .A(N103), .Y(n3506) );
  CLKINVX1 U2597 ( .A(N104), .Y(n3516) );
  CLKINVX1 U2598 ( .A(N105), .Y(n3521) );
  CLKINVX1 U2599 ( .A(N106), .Y(n3526) );
  CLKINVX1 U2600 ( .A(N107), .Y(n3531) );
  CLKINVX1 U2601 ( .A(N180), .Y(n3424) );
  CLKINVX1 U2602 ( .A(N108), .Y(n3536) );
  CLKINVX1 U2603 ( .A(N109), .Y(n3541) );
  CLKINVX1 U2604 ( .A(N110), .Y(n3546) );
  CLKINVX1 U2605 ( .A(N111), .Y(n3551) );
  CLKINVX1 U2606 ( .A(N112), .Y(n3556) );
  CLKINVX1 U2607 ( .A(N113), .Y(n3561) );
  CLKINVX1 U2608 ( .A(N114), .Y(n3408) );
  CLKINVX1 U2609 ( .A(N115), .Y(n3416) );
  CLKINVX1 U2610 ( .A(N116), .Y(n3421) );
  CLKINVX1 U2611 ( .A(N117), .Y(n3426) );
  CLKINVX1 U2612 ( .A(N181), .Y(n3429) );
  CLKINVX1 U2613 ( .A(N118), .Y(n3431) );
  CLKINVX1 U2614 ( .A(N119), .Y(n3436) );
  CLKINVX1 U2615 ( .A(N120), .Y(n3441) );
  CLKINVX1 U2616 ( .A(N121), .Y(n3456) );
  CLKINVX1 U2617 ( .A(N122), .Y(n3511) );
  CLKINVX1 U2618 ( .A(N123), .Y(n3566) );
  CLKINVX1 U2619 ( .A(N124), .Y(n3447) );
  CLKINVX1 U2620 ( .A(N125), .Y(n3452) );
  CLKINVX1 U2621 ( .A(N126), .Y(n3462) );
  CLKINVX1 U2622 ( .A(N127), .Y(n3467) );
  CLKINVX1 U2623 ( .A(N182), .Y(n3434) );
  CLKINVX1 U2624 ( .A(N128), .Y(n3472) );
  CLKINVX1 U2625 ( .A(N129), .Y(n3477) );
  CLKINVX1 U2626 ( .A(N130), .Y(n3482) );
  CLKINVX1 U2627 ( .A(N131), .Y(n3487) );
  CLKINVX1 U2628 ( .A(N132), .Y(n3492) );
  CLKINVX1 U2629 ( .A(N133), .Y(n3497) );
  CLKINVX1 U2630 ( .A(N134), .Y(n3502) );
  CLKINVX1 U2631 ( .A(N135), .Y(n3507) );
  CLKINVX1 U2632 ( .A(N136), .Y(n3517) );
  CLKINVX1 U2633 ( .A(N137), .Y(n3522) );
  CLKINVX1 U2634 ( .A(N183), .Y(n3439) );
  CLKINVX1 U2635 ( .A(N138), .Y(n3527) );
  CLKINVX1 U2636 ( .A(N139), .Y(n3532) );
  CLKINVX1 U2637 ( .A(N140), .Y(n3537) );
  CLKINVX1 U2638 ( .A(N141), .Y(n3542) );
  CLKINVX1 U2639 ( .A(N142), .Y(n3547) );
  CLKINVX1 U2640 ( .A(N143), .Y(n3552) );
  CLKINVX1 U2641 ( .A(N144), .Y(n3557) );
  CLKINVX1 U2642 ( .A(N145), .Y(n3562) );
  CLKINVX1 U2643 ( .A(N146), .Y(n3410) );
  CLKINVX1 U2644 ( .A(N147), .Y(n3417) );
  CLKINVX1 U2645 ( .A(N184), .Y(n3444) );
  CLKINVX1 U2646 ( .A(N148), .Y(n3422) );
  CLKINVX1 U2647 ( .A(N149), .Y(n3427) );
  CLKINVX1 U2648 ( .A(N150), .Y(n3432) );
  CLKINVX1 U2649 ( .A(N151), .Y(n3437) );
  CLKINVX1 U2650 ( .A(N152), .Y(n3442) );
  CLKINVX1 U2651 ( .A(N153), .Y(n3457) );
  CLKINVX1 U2652 ( .A(N154), .Y(n3512) );
  CLKINVX1 U2653 ( .A(N155), .Y(n3567) );
  CLKINVX1 U2654 ( .A(N156), .Y(n3449) );
  CLKINVX1 U2655 ( .A(N157), .Y(n3454) );
  CLKINVX1 U2656 ( .A(N185), .Y(n3459) );
  CLKINVX1 U2657 ( .A(N158), .Y(n3464) );
  CLKINVX1 U2658 ( .A(N159), .Y(n3469) );
  CLKINVX1 U2659 ( .A(N160), .Y(n3474) );
  CLKINVX1 U2660 ( .A(N161), .Y(n3479) );
  CLKINVX1 U2661 ( .A(N162), .Y(n3484) );
  CLKINVX1 U2662 ( .A(N163), .Y(n3489) );
  CLKINVX1 U2663 ( .A(N164), .Y(n3494) );
  CLKINVX1 U2664 ( .A(N165), .Y(n3499) );
  CLKINVX1 U2665 ( .A(N166), .Y(n3504) );
  CLKINVX1 U2666 ( .A(N167), .Y(n3509) );
  CLKINVX1 U2667 ( .A(N186), .Y(n3514) );
  CLKINVX1 U2668 ( .A(N168), .Y(n3519) );
  CLKINVX1 U2669 ( .A(N169), .Y(n3524) );
  CLKINVX1 U2670 ( .A(N170), .Y(n3529) );
  CLKINVX1 U2671 ( .A(N171), .Y(n3534) );
  CLKINVX1 U2672 ( .A(N172), .Y(n3539) );
  CLKINVX1 U2673 ( .A(N173), .Y(n3544) );
  CLKINVX1 U2674 ( .A(N174), .Y(n3549) );
  CLKINVX1 U2675 ( .A(N175), .Y(n3554) );
  CLKINVX1 U2676 ( .A(N60), .Y(n3450) );
  CLKINVX1 U2677 ( .A(N61), .Y(n3455) );
  CLKINVX1 U2678 ( .A(N62), .Y(n3465) );
  CLKINVX1 U2679 ( .A(N63), .Y(n3470) );
  CLKINVX1 U2680 ( .A(N64), .Y(n3475) );
  CLKINVX1 U2681 ( .A(N65), .Y(n3480) );
  CLKINVX1 U2682 ( .A(N66), .Y(n3485) );
  CLKINVX1 U2683 ( .A(N67), .Y(n3490) );
  CLKINVX1 U2684 ( .A(N176), .Y(n3559) );
  CLKINVX1 U2685 ( .A(N68), .Y(n3495) );
  CLKINVX1 U2686 ( .A(N69), .Y(n3500) );
  CLKINVX1 U2687 ( .A(N70), .Y(n3505) );
  CLKINVX1 U2688 ( .A(N71), .Y(n3510) );
  CLKINVX1 U2689 ( .A(N72), .Y(n3520) );
  CLKINVX1 U2690 ( .A(N73), .Y(n3525) );
  CLKINVX1 U2691 ( .A(N74), .Y(n3530) );
  CLKINVX1 U2692 ( .A(N75), .Y(n3535) );
  CLKINVX1 U2693 ( .A(N76), .Y(n3540) );
  CLKINVX1 U2694 ( .A(N77), .Y(n3545) );
  CLKINVX1 U2695 ( .A(N177), .Y(n3564) );
  CLKINVX1 U2696 ( .A(N78), .Y(n3550) );
  CLKINVX1 U2697 ( .A(N79), .Y(n3555) );
  CLKINVX1 U2698 ( .A(N80), .Y(n3560) );
  CLKINVX1 U2699 ( .A(N81), .Y(n3565) );
  CLKINVX1 U2700 ( .A(N82), .Y(n3415) );
  CLKINVX1 U2701 ( .A(N83), .Y(n3420) );
  CLKINVX1 U2702 ( .A(N84), .Y(n3425) );
  CLKINVX1 U2703 ( .A(N85), .Y(n3430) );
  CLKINVX1 U2704 ( .A(N86), .Y(n3435) );
  CLKINVX1 U2705 ( .A(N87), .Y(n3440) );
  CLKINVX1 U2706 ( .A(N187), .Y(n3569) );
  NOR2X1 U2707 ( .A(n413), .B(mem_read), .Y(n3765) );
  NOR3BXL U2708 ( .AN(n3766), .B(n3404), .C(mem_ready), .Y(n6281) );
  NOR2X1 U2709 ( .A(proc_read), .B(proc_write), .Y(n3404) );
  OAI21XL U2710 ( .A0(N34), .A1(n3406), .B0(n3405), .Y(n3766) );
  NAND2BX1 U2711 ( .AN(N33), .B(proc_read), .Y(n3405) );
  CLKINVX1 U2712 ( .A(n3760), .Y(n3406) );
  CLKINVX1 U2713 ( .A(mem_ready), .Y(n3740) );
  NAND4X1 U2714 ( .A(n3768), .B(n3769), .C(n3770), .D(n3771), .Y(n3760) );
  NOR4X1 U2715 ( .A(n3772), .B(n3773), .C(n3774), .D(n3775), .Y(n3771) );
  XOR2X1 U2716 ( .A(proc_addr[25]), .B(N39), .Y(n3775) );
  XOR2X1 U2717 ( .A(proc_addr[23]), .B(N41), .Y(n3774) );
  XOR2X1 U2718 ( .A(proc_addr[24]), .B(N40), .Y(n3773) );
  NAND4X1 U2719 ( .A(n3776), .B(n3777), .C(n3778), .D(n3779), .Y(n3772) );
  XNOR2X1 U2720 ( .A(N35), .B(proc_addr[29]), .Y(n3779) );
  XNOR2X1 U2721 ( .A(N36), .B(proc_addr[28]), .Y(n3778) );
  XNOR2X1 U2722 ( .A(N37), .B(proc_addr[27]), .Y(n3777) );
  XNOR2X1 U2723 ( .A(N38), .B(proc_addr[26]), .Y(n3776) );
  NOR4X1 U2724 ( .A(n3780), .B(n3781), .C(n3782), .D(n3783), .Y(n3770) );
  XOR2X1 U2725 ( .A(proc_addr[19]), .B(N45), .Y(n3783) );
  XOR2X1 U2726 ( .A(proc_addr[17]), .B(N47), .Y(n3782) );
  XOR2X1 U2727 ( .A(proc_addr[18]), .B(N46), .Y(n3781) );
  NAND3X1 U2728 ( .A(n3784), .B(n3785), .C(n3786), .Y(n3780) );
  XNOR2X1 U2729 ( .A(N43), .B(proc_addr[21]), .Y(n3786) );
  XNOR2X1 U2730 ( .A(N44), .B(proc_addr[20]), .Y(n3785) );
  XNOR2X1 U2731 ( .A(N42), .B(proc_addr[22]), .Y(n3784) );
  NOR4X1 U2732 ( .A(n3787), .B(n3788), .C(n3789), .D(n3790), .Y(n3769) );
  XOR2X1 U2733 ( .A(proc_addr[13]), .B(N51), .Y(n3790) );
  XOR2X1 U2734 ( .A(proc_addr[11]), .B(N53), .Y(n3789) );
  XOR2X1 U2735 ( .A(proc_addr[12]), .B(N52), .Y(n3788) );
  NAND3X1 U2736 ( .A(n3791), .B(n3792), .C(n3793), .Y(n3787) );
  XNOR2X1 U2737 ( .A(N49), .B(proc_addr[15]), .Y(n3793) );
  XNOR2X1 U2738 ( .A(N50), .B(proc_addr[14]), .Y(n3792) );
  XNOR2X1 U2739 ( .A(N48), .B(proc_addr[16]), .Y(n3791) );
  NOR4X1 U2740 ( .A(n3794), .B(n3795), .C(n3796), .D(n3797), .Y(n3768) );
  XOR2X1 U2741 ( .A(proc_addr[7]), .B(N57), .Y(n3797) );
  XOR2X1 U2742 ( .A(proc_addr[5]), .B(N59), .Y(n3796) );
  XOR2X1 U2743 ( .A(proc_addr[6]), .B(N58), .Y(n3795) );
  NAND3X1 U2744 ( .A(n3798), .B(n3799), .C(n3800), .Y(n3794) );
  XNOR2X1 U2745 ( .A(N55), .B(proc_addr[9]), .Y(n3800) );
  XNOR2X1 U2746 ( .A(N56), .B(proc_addr[8]), .Y(n3799) );
  XNOR2X1 U2747 ( .A(N54), .B(proc_addr[10]), .Y(n3798) );
  NAND2X1 U2748 ( .A(n3759), .B(n3763), .Y(n3767) );
  NAND2X1 U2749 ( .A(N33), .B(proc_read), .Y(n3763) );
  NAND2X1 U2750 ( .A(proc_write), .B(n3761), .Y(n3759) );
  CLKINVX1 U2751 ( .A(proc_read), .Y(n3761) );
endmodule


module CHIP ( clk, rst_n, mem_read_D, mem_write_D, mem_addr_D, mem_wdata_D, 
        mem_rdata_D, mem_ready_D, mem_read_I, mem_write_I, mem_addr_I, 
        mem_wdata_I, mem_rdata_I, mem_ready_I, DCACHE_addr, DCACHE_wdata, 
        DCACHE_wen );
  output [31:4] mem_addr_D;
  output [127:0] mem_wdata_D;
  input [127:0] mem_rdata_D;
  output [31:4] mem_addr_I;
  output [127:0] mem_wdata_I;
  input [127:0] mem_rdata_I;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input clk, rst_n, mem_ready_D, mem_ready_I;
  output mem_read_D, mem_write_D, mem_read_I, mem_write_I, DCACHE_wen;
  wire   n7, n8, n9, n10, n11, ICACHE_stall, DCACHE_ren, DCACHE_stall, n1;
  wire   [29:0] ICACHE_addr;
  wire   [31:0] ICACHE_wdata;
  wire   [31:0] ICACHE_rdata;
  wire   [31:0] DCACHE_rdata;

  MIPS_Pipeline i_MIPS ( .clk(clk), .rst_n(rst_n), .ICACHE_addr(ICACHE_addr), 
        .ICACHE_stall(ICACHE_stall), .ICACHE_rdata(ICACHE_rdata), .DCACHE_ren(
        DCACHE_ren), .DCACHE_wen(DCACHE_wen), .DCACHE_addr({DCACHE_addr[29:5], 
        n9, n10, n11, DCACHE_addr[1:0]}), .DCACHE_wdata(DCACHE_wdata), 
        .DCACHE_stall(DCACHE_stall), .DCACHE_rdata(DCACHE_rdata) );
  cache_0 D_cache ( .clk(clk), .proc_reset(n1), .proc_read(DCACHE_ren), 
        .proc_write(DCACHE_wen), .proc_addr(DCACHE_addr), .proc_wdata(
        DCACHE_wdata), .proc_stall(DCACHE_stall), .proc_rdata(DCACHE_rdata), 
        .mem_read(mem_read_D), .mem_write(n7), .mem_addr(mem_addr_D), 
        .mem_rdata(mem_rdata_D), .mem_wdata(mem_wdata_D), .mem_ready(
        mem_ready_D) );
  cache_1 I_cache ( .clk(clk), .proc_reset(n1), .proc_read(1'b1), .proc_write(
        1'b0), .proc_addr(ICACHE_addr), .proc_wdata({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .proc_stall(ICACHE_stall), .proc_rdata(
        ICACHE_rdata), .mem_read(mem_read_I), .mem_write(n8), .mem_addr(
        mem_addr_I), .mem_rdata(mem_rdata_I), .mem_wdata(mem_wdata_I), 
        .mem_ready(mem_ready_I) );
  BUFX12 U2 ( .A(n10), .Y(DCACHE_addr[3]) );
  BUFX12 U3 ( .A(n9), .Y(DCACHE_addr[4]) );
  BUFX12 U4 ( .A(n8), .Y(mem_write_I) );
  BUFX12 U5 ( .A(n7), .Y(mem_write_D) );
  BUFX16 U6 ( .A(n11), .Y(DCACHE_addr[2]) );
  CLKINVX1 U7 ( .A(rst_n), .Y(n1) );
endmodule

