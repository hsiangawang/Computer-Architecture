module settmine (mine_number,set_ready);

input reg [3:0] mine_number;
output reg  set_ready;



